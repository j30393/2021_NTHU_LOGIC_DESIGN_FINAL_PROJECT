module ball_display(
    input [15:0]pos,
    output reg white
);



always@(*)begin

    if(pos==264||
        pos==265||pos==313||pos==314||pos==315||pos==362||pos==363||
        pos==364||pos==365||pos==377||pos==378||pos==412||pos==413||
        pos==414||pos==415||pos==426||pos==427||pos==428||pos==462||
        pos==463||pos==464||pos==465||pos==475||pos==476||pos==477||
        pos==478||pos==511||pos==512||pos==513||pos==514||pos==524||
        pos==525||pos==526||pos==527||pos==528||pos==561||pos==562||
        pos==563||pos==564||pos==566||pos==567||pos==568||pos==569||
        pos==570||pos==571||pos==572||pos==573||pos==574||pos==575||
        pos==576||pos==577||pos==578||pos==611||pos==612||pos==613||
        pos==614||pos==615||pos==616||pos==617||pos==618||pos==619||
        pos==620||pos==621||pos==622||pos==623||pos==624||pos==625||
        pos==626||pos==627||pos==661||pos==662||pos==663||pos==664||
        pos==665||pos==666||pos==667||pos==668||pos==669||pos==670||
        pos==671||pos==672||pos==673||pos==674||pos==675||pos==676||
        pos==677||pos==711||pos==712||pos==713||pos==714||pos==715||
        pos==716||pos==717||pos==718||pos==719||pos==720||pos==721||
        pos==722||pos==723||pos==724||pos==725||pos==726||pos==727||
        pos==761||pos==762||pos==763||pos==764||pos==765||pos==766||
        pos==767||pos==768||pos==769||pos==770||pos==771||pos==772||
        pos==773||pos==774||pos==775||pos==776||pos==777||pos==778||
        pos==811||pos==812||pos==813||pos==814||pos==815||pos==816||
        pos==817||pos==818||pos==819||pos==820||pos==821||pos==822||
        pos==823||pos==824||pos==825||pos==826||pos==827||pos==828||
        pos==829||pos==860||pos==861||pos==862||pos==863||pos==864||
        pos==865||pos==866||pos==867||pos==868||pos==869||pos==870||
        pos==871||pos==872||pos==873||pos==874||pos==875||pos==876||
        pos==877||pos==878||pos==879||pos==910||pos==911||pos==912||
        pos==913||pos==914||pos==915||pos==916||pos==917||pos==918||
        pos==919||pos==920||pos==921||pos==922||pos==923||pos==924||
        pos==925||pos==926||pos==927||pos==928||pos==929||pos==930||
        pos==959||pos==960||pos==961||pos==962||pos==963||pos==964||
        pos==965||pos==966||pos==967||pos==968||pos==969||pos==970||
        pos==971||pos==972||pos==973||pos==974||pos==975||pos==976||
        pos==977||pos==978||pos==979||pos==980||pos==1009||pos==1010||
        pos==1011||pos==1012||pos==1013||pos==1014||pos==1015||pos==1016||
        pos==1017||pos==1018||pos==1019||pos==1020||pos==1021||pos==1022||
        pos==1023||pos==1024||pos==1025||pos==1026||pos==1027||pos==1028||
        pos==1029||pos==1030||pos==1031||pos==1058||pos==1059||pos==1060||
        pos==1061||pos==1062||pos==1063||pos==1064||pos==1065||pos==1066||
        pos==1067||pos==1068||pos==1069||pos==1070||pos==1071||pos==1072||
        pos==1073||pos==1074||pos==1075||pos==1076||pos==1077||pos==1078||
        pos==1079||pos==1080||pos==1081||pos==1108||pos==1109||pos==1110||
        pos==1111||pos==1112||pos==1113||pos==1114||pos==1115||pos==1116||
        pos==1117||pos==1118||pos==1119||pos==1120||pos==1121||pos==1122||
        pos==1123||pos==1124||pos==1125||pos==1126||pos==1127||pos==1128||
        pos==1129||pos==1130||pos==1131||pos==1157||pos==1158||pos==1159||
        pos==1160||pos==1161||pos==1162||pos==1163||pos==1164||pos==1165||
        pos==1166||pos==1167||pos==1168||pos==1169||pos==1170||pos==1171||
        pos==1172||pos==1173||pos==1174||pos==1175||pos==1176||pos==1177||
        pos==1178||pos==1179||pos==1180||pos==1181||pos==1182||pos==1207||
        pos==1208||pos==1209||pos==1210||pos==1211||pos==1212||pos==1213||
        pos==1214||pos==1215||pos==1216||pos==1217||pos==1218||pos==1219||
        pos==1220||pos==1221||pos==1222||pos==1223||pos==1224||pos==1225||
        pos==1226||pos==1227||pos==1228||pos==1229||pos==1230||pos==1231||
        pos==1232||pos==1257||pos==1258||pos==1259||pos==1260||pos==1261||
        pos==1262||pos==1263||pos==1264||pos==1265||pos==1266||pos==1267||
        pos==1268||pos==1269||pos==1270||pos==1271||pos==1272||pos==1273||
        pos==1274||pos==1275||pos==1276||pos==1277||pos==1278||pos==1279||
        pos==1280||pos==1281||pos==1282||pos==1292||pos==1293||pos==1294||
        pos==1295||pos==1307||pos==1308||pos==1309||pos==1310||pos==1311||
        pos==1312||pos==1313||pos==1314||pos==1315||pos==1316||pos==1317||
        pos==1318||pos==1319||pos==1320||pos==1321||pos==1322||pos==1323||
        pos==1324||pos==1325||pos==1326||pos==1327||pos==1328||pos==1329||
        pos==1330||pos==1331||pos==1332||pos==1339||pos==1340||pos==1341||
        pos==1342||pos==1343||pos==1344||pos==1345||pos==1346||pos==1357||
        pos==1358||pos==1359||pos==1360||pos==1361||pos==1362||pos==1363||
        pos==1364||pos==1365||pos==1366||pos==1367||pos==1368||pos==1369||
        pos==1370||pos==1371||pos==1372||pos==1373||pos==1374||pos==1375||
        pos==1376||pos==1377||pos==1378||pos==1379||pos==1380||pos==1381||
        pos==1382||pos==1386||pos==1387||pos==1388||pos==1389||pos==1390||
        pos==1391||pos==1392||pos==1393||pos==1394||pos==1395||pos==1396||
        pos==1407||pos==1408||pos==1409||pos==1410||pos==1411||pos==1412||
        pos==1413||pos==1414||pos==1415||pos==1416||pos==1417||pos==1418||
        pos==1419||pos==1420||pos==1421||pos==1422||pos==1423||pos==1424||
        pos==1425||pos==1426||pos==1427||pos==1428||pos==1429||pos==1430||
        pos==1431||pos==1432||pos==1436||pos==1437||pos==1438||pos==1439||
        pos==1440||pos==1441||pos==1442||pos==1443||pos==1444||pos==1445||
        pos==1446||pos==1457||pos==1458||pos==1459||pos==1460||pos==1461||
        pos==1462||pos==1463||pos==1464||pos==1465||pos==1466||pos==1467||
        pos==1468||pos==1469||pos==1470||pos==1471||pos==1472||pos==1473||
        pos==1474||pos==1475||pos==1476||pos==1477||pos==1478||pos==1479||
        pos==1480||pos==1481||pos==1482||pos==1486||pos==1487||pos==1488||
        pos==1489||pos==1490||pos==1491||pos==1492||pos==1493||pos==1494||
        pos==1495||pos==1506||pos==1507||pos==1508||pos==1509||pos==1510||
        pos==1511||pos==1512||pos==1513||pos==1514||pos==1515||pos==1516||
        pos==1517||pos==1518||pos==1519||pos==1520||pos==1521||pos==1522||
        pos==1523||pos==1524||pos==1525||pos==1526||pos==1527||pos==1528||
        pos==1529||pos==1530||pos==1531||pos==1532||pos==1536||pos==1537||
        pos==1538||pos==1539||pos==1540||pos==1541||pos==1542||pos==1543||
        pos==1544||pos==1545||pos==1556||pos==1557||pos==1558||pos==1559||
        pos==1560||pos==1561||pos==1562||pos==1563||pos==1564||pos==1565||
        pos==1566||pos==1567||pos==1568||pos==1569||pos==1570||pos==1571||
        pos==1572||pos==1573||pos==1574||pos==1575||pos==1576||pos==1577||
        pos==1578||pos==1579||pos==1580||pos==1581||pos==1582||pos==1585||
        pos==1586||pos==1587||pos==1588||pos==1589||pos==1590||pos==1591||
        pos==1592||pos==1593||pos==1594||pos==1595||pos==1606||pos==1607||
        pos==1608||pos==1609||pos==1610||pos==1611||pos==1612||pos==1613||
        pos==1614||pos==1615||pos==1616||pos==1617||pos==1618||pos==1619||
        pos==1620||pos==1621||pos==1622||pos==1623||pos==1624||pos==1625||
        pos==1626||pos==1627||pos==1628||pos==1629||pos==1630||pos==1631||
        pos==1632||pos==1633||pos==1634||pos==1635||pos==1636||pos==1637||
        pos==1638||pos==1639||pos==1640||pos==1641||pos==1642||pos==1643||
        pos==1644||pos==1645||pos==1657||pos==1658||pos==1659||pos==1660||
        pos==1661||pos==1662||pos==1663||pos==1664||pos==1665||pos==1666||
        pos==1667||pos==1668||pos==1669||pos==1670||pos==1671||pos==1672||
        pos==1673||pos==1674||pos==1675||pos==1676||pos==1677||pos==1678||
        pos==1679||pos==1680||pos==1681||pos==1682||pos==1683||pos==1684||
        pos==1685||pos==1686||pos==1687||pos==1688||pos==1689||pos==1690||
        pos==1691||pos==1692||pos==1693||pos==1694||pos==1695||pos==1707||
        pos==1708||pos==1709||pos==1710||pos==1711||pos==1712||pos==1713||
        pos==1714||pos==1715||pos==1716||pos==1717||pos==1718||pos==1719||
        pos==1720||pos==1721||pos==1722||pos==1723||pos==1724||pos==1725||
        pos==1726||pos==1727||pos==1728||pos==1729||pos==1730||pos==1731||
        pos==1732||pos==1733||pos==1734||pos==1735||pos==1736||pos==1737||
        pos==1738||pos==1739||pos==1740||pos==1741||pos==1742||pos==1743||
        pos==1744||pos==1757||pos==1758||pos==1759||pos==1760||pos==1761||
        pos==1762||pos==1763||pos==1764||pos==1765||pos==1766||pos==1767||
        pos==1768||pos==1769||pos==1770||pos==1771||pos==1772||pos==1773||
        pos==1774||pos==1775||pos==1776||pos==1777||pos==1778||pos==1779||
        pos==1780||pos==1781||pos==1782||pos==1783||pos==1784||pos==1785||
        pos==1790||pos==1791||pos==1792||pos==1793||pos==1794||pos==1807||
        pos==1808||pos==1809||pos==1810||pos==1811||pos==1812||pos==1813||
        pos==1814||pos==1815||pos==1816||pos==1817||pos==1818||pos==1819||
        pos==1820||pos==1821||pos==1822||pos==1823||pos==1824||pos==1825||
        pos==1826||pos==1827||pos==1828||pos==1829||pos==1830||pos==1831||
        pos==1833||pos==1834||pos==1835||pos==1842||pos==1843||pos==1844||
        pos==1858||pos==1859||pos==1860||pos==1861||pos==1862||pos==1863||
        pos==1864||pos==1865||pos==1866||pos==1867||pos==1868||pos==1869||
        pos==1870||pos==1871||pos==1872||pos==1873||pos==1874||pos==1875||
        pos==1876||pos==1877||pos==1878||pos==1879||pos==1880||pos==1881||
        pos==1893||pos==1908||pos==1909||pos==1910||pos==1911||pos==1912||
        pos==1913||pos==1914||pos==1915||pos==1916||pos==1917||pos==1918||
        pos==1919||pos==1920||pos==1921||pos==1922||pos==1923||pos==1924||
        pos==1925||pos==1926||pos==1927||pos==1928||pos==1929||pos==1930||
        pos==1958||pos==1959||pos==1960||pos==1961||pos==1962||pos==1963||
        pos==1964||pos==1965||pos==1966||pos==1967||pos==1968||pos==1969||
        pos==1970||pos==1971||pos==1972||pos==1973||pos==1974||pos==1975||
        pos==1976||pos==1977||pos==1978||pos==1979||pos==2008||pos==2009||
        pos==2010||pos==2011||pos==2012||pos==2013||pos==2014||pos==2015||
        pos==2016||pos==2017||pos==2018||pos==2019||pos==2020||pos==2021||
        pos==2022||pos==2023||pos==2024||pos==2025||pos==2026||pos==2027||
        pos==2028||pos==2029||pos==2059||pos==2060||pos==2061||pos==2062||
        pos==2063||pos==2064||pos==2065||pos==2066||pos==2067||pos==2068||
        pos==2069||pos==2070||pos==2071||pos==2072||pos==2073||pos==2074||
        pos==2075||pos==2076||pos==2077||pos==2078||pos==2079||pos==2109||
        pos==2110||pos==2111||pos==2112||pos==2113||pos==2114||pos==2115||
        pos==2116||pos==2117||pos==2118||pos==2119||pos==2120||pos==2121||
        pos==2122||pos==2123||pos==2124||pos==2125||pos==2126||pos==2127||
        pos==2128||pos==2129||pos==2160||pos==2161||pos==2162||pos==2163||
        pos==2164||pos==2165||pos==2166||pos==2167||pos==2168||pos==2169||
        pos==2170||pos==2171||pos==2172||pos==2173||pos==2174||pos==2175||
        pos==2176||pos==2177||pos==2179||pos==2211||pos==2212||pos==2213||
        pos==2214||pos==2215||pos==2216||pos==2217||pos==2218||pos==2219||
        pos==2220||pos==2221||pos==2222||pos==2223||pos==2224||pos==2225||
        pos==2226||pos==2262||pos==2263||pos==2264||pos==2265||pos==2266||
        pos==2267||pos==2268||pos==2269||pos==2270||pos==2271||pos==2272||
        pos==2273||pos==2274||pos==2313||pos==2314||pos==2315||pos==2316||
        pos==2317||pos==2318||pos==2319||pos==2320||pos==2321||pos==2322||
        pos==2323||pos==2324||pos==2366||pos==2367||pos==2368||pos==2369) white=0;
    else white=1;

end

endmodule