`define lllc  32'd32  // C1
`define llc  32'd65  // C2
`define llf  32'd87   // F2
`define llg  32'd98   // G2
`define lla  32'd110   // A2
`define llb  32'd123   // B2
`define lc  32'd131   // C3
`define ld  32'd147   // C3
`define le  32'd165   // C3
`define lf  32'd174   // F3
`define lg  32'd196  // G3
`define la  32'd220   // C3
`define lsa   32'd233   // #A3
`define lb  32'd247   // C3
`define c   32'd262   // C4
`define d   32'd294   // D4
`define e   32'd330   // E4
`define f   32'd349   // F4
`define sf   32'd370   // #F4
`define g   32'd392   // G4
`define a   32'd440   // A4
`define sa   32'd466   // #A4
`define b   32'd494   // B4
`define hc   32'd524   // C4
`define hd   32'd588   // D4
`define he   32'd660   // E4
`define hf   32'd698   // F4
`define hg   32'd784   // G4
`define ha   32'd880   // A4
`define hb   32'd988   // B4


`define sil   32'd50000000 // slience

module music_example (
	input [11:0] ibeatNum,
    input en,
	output reg [31:0] toneL,
    output reg [31:0] toneR
);

always @(*) begin
    if(en) begin
        case(ibeatNum)
                12'd0: toneR = `g;
                12'd1: toneR = `g;
                12'd2: toneR = `g;
                12'd3: toneR = `g;
                12'd4: toneR = `sf;
                12'd5: toneR = `sf;
                12'd6: toneR = `sf;
                12'd7: toneR = `sf;
                12'd8: toneR = `g;
                12'd9: toneR = `g;
                12'd10: toneR = `g;
                12'd11: toneR = `g;
                12'd12: toneR = `a;
                12'd13: toneR = `a;
                12'd14: toneR = `a;
                12'd15: toneR = `a;
                12'd16: toneR = `g;
                12'd17: toneR = `g;
                12'd18: toneR = `g;
                12'd19: toneR = `g;
                12'd20: toneR = `g;
                12'd21: toneR = `g;
                12'd22: toneR = `g;
                12'd23: toneR = `g;
                12'd24: toneR = `g;
                12'd25: toneR = `g;
                12'd26: toneR = `g;
                12'd27: toneR = `g;
                12'd28: toneR = `sil;
                12'd29: toneR = `sil;
                12'd30: toneR = `sil;
                12'd31: toneR = `sil;
                12'd32: toneR = `g;
                12'd33: toneR = `g;
                12'd34: toneR = `g;
                12'd35: toneR = `g;
                12'd36: toneR = `sf;
                12'd37: toneR = `sf;
                12'd38: toneR = `sf;
                12'd39: toneR = `sf;
                12'd40: toneR = `g;
                12'd41: toneR = `g;
                12'd42: toneR = `g;
                12'd43: toneR = `g;
                12'd44: toneR = `a;
                12'd45: toneR = `a;
                12'd46: toneR = `a;
                12'd47: toneR = `a;
                12'd48: toneR = `g;
                12'd49: toneR = `g;
                12'd50: toneR = `g;
                12'd51: toneR = `g;
                12'd52: toneR = `g;
                12'd53: toneR = `g;
                12'd54: toneR = `g;
                12'd55: toneR = `g;
                12'd56: toneR = `g;
                12'd57: toneR = `g;
                12'd58: toneR = `g;
                12'd59: toneR = `g;
                12'd60: toneR = `sil;
                12'd61: toneR = `sil;
                12'd62: toneR = `sil;
                12'd63: toneR = `sil;
                12'd64: toneR = `g;
                12'd65: toneR = `g;
                12'd66: toneR = `g;
                12'd67: toneR = `sil;
                12'd68: toneR = `g;
                12'd69: toneR = `g;
                12'd70: toneR = `g;
                12'd71: toneR = `sil;
                12'd72: toneR = `g;
                12'd73: toneR = `g;
                12'd74: toneR = `g;
                12'd75: toneR = `g;
                12'd76: toneR = `g;
                12'd77: toneR = `g;
                12'd78: toneR = `g;
                12'd79: toneR = `g;
                12'd80: toneR = `a;
                12'd81: toneR = `a;
                12'd82: toneR = `a;
                12'd83: toneR = `a;
                12'd84: toneR = `a;
                12'd85: toneR = `a;
                12'd86: toneR = `a;
                12'd87: toneR = `a;
                12'd88: toneR = `sa;
                12'd89: toneR = `sa;
                12'd90: toneR = `sa;
                12'd91: toneR = `sa;
                12'd92: toneR = `sa;
                12'd93: toneR = `sa;
                12'd94: toneR = `sa;
                12'd95: toneR = `sa;
                12'd96: toneR = `b;
                12'd97: toneR = `b;
                12'd98: toneR = `b;
                12'd99: toneR = `b;
                12'd100: toneR = `b;
                12'd101: toneR = `b;
                12'd102: toneR = `b;
                12'd103: toneR = `b;
                12'd104: toneR = `g;
                12'd105: toneR = `g;
                12'd106: toneR = `g;
                12'd107: toneR = `g;
                12'd108: toneR = `g;
                12'd109: toneR = `g;
                12'd110: toneR = `g;
                12'd111: toneR = `g;
                12'd112: toneR = `a;
                12'd113: toneR = `a;
                12'd114: toneR = `a;
                12'd115: toneR = `a;
                12'd116: toneR = `a;
                12'd117: toneR = `a;
                12'd118: toneR = `a;
                12'd119: toneR = `a;
                12'd120: toneR = `b;
                12'd121: toneR = `b;
                12'd122: toneR = `b;
                12'd123: toneR = `b;
                12'd124: toneR = `b;
                12'd125: toneR = `b;
                12'd126: toneR = `b;
                12'd127: toneR = `b;
                12'd128: toneR = `hc;
                12'd129: toneR = `hc;
                12'd130: toneR = `hc;
                12'd131: toneR = `hc;
                12'd132: toneR = `hc;
                12'd133: toneR = `hc;
                12'd134: toneR = `hc;
                12'd135: toneR = `hc;
                12'd136: toneR = `b;
                12'd137: toneR = `b;
                12'd138: toneR = `b;
                12'd139: toneR = `b;
                12'd140: toneR = `b;
                12'd141: toneR = `b;
                12'd142: toneR = `b;
                12'd143: toneR = `b;
                12'd144: toneR = `hc;
                12'd145: toneR = `hc;
                12'd146: toneR = `hc;
                12'd147: toneR = `hc;
                12'd148: toneR = `hc;
                12'd149: toneR = `hc;
                12'd150: toneR = `hc;
                12'd151: toneR = `hc;
                12'd152: toneR = `b;
                12'd153: toneR = `b;
                12'd154: toneR = `b;
                12'd155: toneR = `b;
                12'd156: toneR = `hc;
                12'd157: toneR = `hc;
                12'd158: toneR = `hc;
                12'd159: toneR = `hc;
                12'd160: toneR = `sil;
                12'd161: toneR = `sil;
                12'd162: toneR = `sil;
                12'd163: toneR = `sil;
                12'd164: toneR = `sil;
                12'd165: toneR = `sil;
                12'd166: toneR = `sil;
                12'd167: toneR = `sil;
                12'd168: toneR = `b;
                12'd169: toneR = `b;
                12'd170: toneR = `b;
                12'd171: toneR = `b;
                12'd172: toneR = `b;
                12'd173: toneR = `b;
                12'd174: toneR = `b;
                12'd175: toneR = `b;
                12'd176: toneR = `hc;
                12'd177: toneR = `hc;
                12'd178: toneR = `hc;
                12'd179: toneR = `hc;
                12'd180: toneR = `hc;
                12'd181: toneR = `hc;
                12'd182: toneR = `hc;
                12'd183: toneR = `hc;
                12'd184: toneR = `b;
                12'd185: toneR = `b;
                12'd186: toneR = `b;
                12'd187: toneR = `b;
                12'd188: toneR = `b;
                12'd189: toneR = `b;
                12'd190: toneR = `b;
                12'd191: toneR = `b;
                12'd192: toneR = `a;
                12'd193: toneR = `a;
                12'd194: toneR = `a;
                12'd195: toneR = `a;
                12'd196: toneR = `a;
                12'd197: toneR = `a;
                12'd198: toneR = `a;
                12'd199: toneR = `a;
                12'd200: toneR = `g;
                12'd201: toneR = `g;
                12'd202: toneR = `g;
                12'd203: toneR = `g;
                12'd204: toneR = `g;
                12'd205: toneR = `g;
                12'd206: toneR = `g;
                12'd207: toneR = `g;
                12'd208: toneR = `a;
                12'd209: toneR = `a;
                12'd210: toneR = `a;
                12'd211: toneR = `a;
                12'd212: toneR = `a;
                12'd213: toneR = `a;
                12'd214: toneR = `a;
                12'd215: toneR = `a;
                12'd216: toneR = `g;
                12'd217: toneR = `g;
                12'd218: toneR = `g;
                12'd219: toneR = `g;
                12'd220: toneR = `a;
                12'd221: toneR = `a;
                12'd222: toneR = `a;
                12'd223: toneR = `a;
                12'd224: toneR = `sil;
                12'd225: toneR = `sil;
                12'd226: toneR = `sil;
                12'd227: toneR = `sil;
                12'd228: toneR = `sil;
                12'd229: toneR = `sil;
                12'd230: toneR = `sil;
                12'd231: toneR = `sil;
                12'd232: toneR = `g;
                12'd233: toneR = `g;
                12'd234: toneR = `g;
                12'd235: toneR = `g;
                12'd236: toneR = `g;
                12'd237: toneR = `g;
                12'd238: toneR = `g;
                12'd239: toneR = `g;
                12'd240: toneR = `a;
                12'd241: toneR = `a;
                12'd242: toneR = `a;
                12'd243: toneR = `a;
                12'd244: toneR = `a;
                12'd245: toneR = `a;
                12'd246: toneR = `a;
                12'd247: toneR = `a;
                12'd248: toneR = `b;
                12'd249: toneR = `b;
                12'd250: toneR = `b;
                12'd251: toneR = `b;
                12'd252: toneR = `b;
                12'd253: toneR = `b;
                12'd254: toneR = `b;
                12'd255: toneR = `b;
                12'd256: toneR = `hc;
                12'd257: toneR = `hc;
                12'd258: toneR = `hc;
                12'd259: toneR = `hc;
                12'd260: toneR = `hc;
                12'd261: toneR = `hc;
                12'd262: toneR = `hc;
                12'd263: toneR = `hc;
                12'd264: toneR = `b;
                12'd265: toneR = `b;
                12'd266: toneR = `b;
                12'd267: toneR = `b;
                12'd268: toneR = `b;
                12'd269: toneR = `b;
                12'd270: toneR = `b;
                12'd271: toneR = `b;
                12'd272: toneR = `hc;
                12'd273: toneR = `hc;
                12'd274: toneR = `hc;
                12'd275: toneR = `hc;
                12'd276: toneR = `hc;
                12'd277: toneR = `hc;
                12'd278: toneR = `hc;
                12'd279: toneR = `hc;
                12'd280: toneR = `b;
                12'd281: toneR = `b;
                12'd282: toneR = `b;
                12'd283: toneR = `b;
                12'd284: toneR = `hc;
                12'd285: toneR = `hc;
                12'd286: toneR = `hc;
                12'd287: toneR = `hc;
                12'd288: toneR = `sil;
                12'd289: toneR = `sil;
                12'd290: toneR = `sil;
                12'd291: toneR = `sil;
                12'd292: toneR = `sil;
                12'd293: toneR = `sil;
                12'd294: toneR = `sil;
                12'd295: toneR = `sil;
                12'd296: toneR = `b;
                12'd297: toneR = `b;
                12'd298: toneR = `b;
                12'd299: toneR = `b;
                12'd300: toneR = `b;
                12'd301: toneR = `b;
                12'd302: toneR = `b;
                12'd303: toneR = `b;
                12'd304: toneR = `hc;
                12'd305: toneR = `hc;
                12'd306: toneR = `hc;
                12'd307: toneR = `hc;
                12'd308: toneR = `hc;
                12'd309: toneR = `hc;
                12'd310: toneR = `hc;
                12'd311: toneR = `hc;
                12'd312: toneR = `b;
                12'd313: toneR = `b;
                12'd314: toneR = `b;
                12'd315: toneR = `b;
                12'd316: toneR = `b;
                12'd317: toneR = `b;
                12'd318: toneR = `b;
                12'd319: toneR = `b;
                12'd320: toneR = `a;
                12'd321: toneR = `a;
                12'd322: toneR = `a;
                12'd323: toneR = `a;
                12'd324: toneR = `a;
                12'd325: toneR = `a;
                12'd326: toneR = `a;
                12'd327: toneR = `a;
                12'd328: toneR = `g;
                12'd329: toneR = `g;
                12'd330: toneR = `g;
                12'd331: toneR = `g;
                12'd332: toneR = `g;
                12'd333: toneR = `g;
                12'd334: toneR = `g;
                12'd335: toneR = `g;
                12'd336: toneR = `a;
                12'd337: toneR = `a;
                12'd338: toneR = `a;
                12'd339: toneR = `a;
                12'd340: toneR = `a;
                12'd341: toneR = `a;
                12'd342: toneR = `a;
                12'd343: toneR = `a;
                12'd344: toneR = `g;
                12'd345: toneR = `g;
                12'd346: toneR = `g;
                12'd347: toneR = `g;
                12'd348: toneR = `a;
                12'd349: toneR = `a;
                12'd350: toneR = `a;
                12'd351: toneR = `a;
                12'd352: toneR = `sil;
                12'd353: toneR = `sil;
                12'd354: toneR = `sil;
                12'd355: toneR = `sil;
                12'd356: toneR = `sil;
                12'd357: toneR = `sil;
                12'd358: toneR = `sil;
                12'd359: toneR = `sil;
                12'd360: toneR = `g;
                12'd361: toneR = `g;
                12'd362: toneR = `g;
                12'd363: toneR = `g;
                12'd364: toneR = `g;
                12'd365: toneR = `g;
                12'd366: toneR = `g;
                12'd367: toneR = `g;
                12'd368: toneR = `a;
                12'd369: toneR = `a;
                12'd370: toneR = `a;
                12'd371: toneR = `a;
                12'd372: toneR = `a;
                12'd373: toneR = `a;
                12'd374: toneR = `a;
                12'd375: toneR = `a;
                12'd376: toneR = `b;
                12'd377: toneR = `b;
                12'd378: toneR = `b;
                12'd379: toneR = `b;
                12'd380: toneR = `b;
                12'd381: toneR = `b;
                12'd382: toneR = `b;
                12'd383: toneR = `b;
                12'd384: toneR = `hc;
                12'd385: toneR = `hc;
                12'd386: toneR = `hc;
                12'd387: toneR = `hc;
                12'd388: toneR = `hc;
                12'd389: toneR = `hc;
                12'd390: toneR = `hc;
                12'd391: toneR = `hc;
                12'd392: toneR = `b;
                12'd393: toneR = `b;
                12'd394: toneR = `b;
                12'd395: toneR = `b;
                12'd396: toneR = `b;
                12'd397: toneR = `b;
                12'd398: toneR = `b;
                12'd399: toneR = `b;
                12'd400: toneR = `hc;
                12'd401: toneR = `hc;
                12'd402: toneR = `hc;
                12'd403: toneR = `hc;
                12'd404: toneR = `hc;
                12'd405: toneR = `hc;
                12'd406: toneR = `hc;
                12'd407: toneR = `hc;
                12'd408: toneR = `b;
                12'd409: toneR = `b;
                12'd410: toneR = `b;
                12'd411: toneR = `b;
                12'd412: toneR = `hc;
                12'd413: toneR = `hc;
                12'd414: toneR = `hc;
                12'd415: toneR = `hc;
                12'd416: toneR = `sil;
                12'd417: toneR = `sil;
                12'd418: toneR = `sil;
                12'd419: toneR = `sil;
                12'd420: toneR = `sil;
                12'd421: toneR = `sil;
                12'd422: toneR = `sil;
                12'd423: toneR = `sil;
                12'd424: toneR = `b;
                12'd425: toneR = `b;
                12'd426: toneR = `b;
                12'd427: toneR = `b;
                12'd428: toneR = `b;
                12'd429: toneR = `b;
                12'd430: toneR = `b;
                12'd431: toneR = `b;
                12'd432: toneR = `hc;
                12'd433: toneR = `hc;
                12'd434: toneR = `hc;
                12'd435: toneR = `hc;
                12'd436: toneR = `hc;
                12'd437: toneR = `hc;
                12'd438: toneR = `hc;
                12'd439: toneR = `hc;
                12'd440: toneR = `b;
                12'd441: toneR = `b;
                12'd442: toneR = `b;
                12'd443: toneR = `b;
                12'd444: toneR = `b;
                12'd445: toneR = `b;
                12'd446: toneR = `b;
                12'd447: toneR = `b;
                12'd448: toneR = `a;
                12'd449: toneR = `a;
                12'd450: toneR = `a;
                12'd451: toneR = `a;
                12'd452: toneR = `a;
                12'd453: toneR = `a;
                12'd454: toneR = `a;
                12'd455: toneR = `a;
                12'd456: toneR = `g;
                12'd457: toneR = `g;
                12'd458: toneR = `g;
                12'd459: toneR = `g;
                12'd460: toneR = `g;
                12'd461: toneR = `g;
                12'd462: toneR = `g;
                12'd463: toneR = `g;
                12'd464: toneR = `a;
                12'd465: toneR = `a;
                12'd466: toneR = `a;
                12'd467: toneR = `a;
                12'd468: toneR = `a;
                12'd469: toneR = `a;
                12'd470: toneR = `a;
                12'd471: toneR = `a;
                12'd472: toneR = `g;
                12'd473: toneR = `g;
                12'd474: toneR = `g;
                12'd475: toneR = `g;
                12'd476: toneR = `a;
                12'd477: toneR = `a;
                12'd478: toneR = `a;
                12'd479: toneR = `a;
                12'd480: toneR = `sil;
                12'd481: toneR = `sil;
                12'd482: toneR = `sil;
                12'd483: toneR = `sil;
                12'd484: toneR = `sil;
                12'd485: toneR = `sil;
                12'd486: toneR = `sil;
                12'd487: toneR = `sil;
                12'd488: toneR = `g;
                12'd489: toneR = `g;
                12'd490: toneR = `g;
                12'd491: toneR = `g;
                12'd492: toneR = `g;
                12'd493: toneR = `g;
                12'd494: toneR = `g;
                12'd495: toneR = `g;
                12'd496: toneR = `a;
                12'd497: toneR = `a;
                12'd498: toneR = `a;
                12'd499: toneR = `a;
                12'd500: toneR = `a;
                12'd501: toneR = `a;
                12'd502: toneR = `a;
                12'd503: toneR = `a;
                12'd504: toneR = `b;
                12'd505: toneR = `b;
                12'd506: toneR = `b;
                12'd507: toneR = `b;
                12'd508: toneR = `b;
                12'd509: toneR = `b;
                12'd510: toneR = `b;
                12'd511: toneR = `b;
                12'd512: toneR = `e;
                12'd513: toneR = `e;
                12'd514: toneR = `e;
                12'd515: toneR = `e;
                12'd516: toneR = `e;
                12'd517: toneR = `e;
                12'd518: toneR = `e;
                12'd519: toneR = `sil;
                12'd520: toneR = `e;
                12'd521: toneR = `e;
                12'd522: toneR = `e;
                12'd523: toneR = `e;
                12'd524: toneR = `e;
                12'd525: toneR = `e;
                12'd526: toneR = `e;
                12'd527: toneR = `e;
                12'd528: toneR = `f;
                12'd529: toneR = `f;
                12'd530: toneR = `f;
                12'd531: toneR = `f;
                12'd532: toneR = `f;
                12'd533: toneR = `f;
                12'd534: toneR = `f;
                12'd535: toneR = `f;
                12'd536: toneR = `g;
                12'd537: toneR = `g;
                12'd538: toneR = `g;
                12'd539: toneR = `g;
                12'd540: toneR = `g;
                12'd541: toneR = `g;
                12'd542: toneR = `g;
                12'd543: toneR = `g;
                12'd544: toneR = `c;
                12'd545: toneR = `c;
                12'd546: toneR = `c;
                12'd547: toneR = `c;
                12'd548: toneR = `c;
                12'd549: toneR = `c;
                12'd550: toneR = `c;
                12'd551: toneR = `c;
                12'd552: toneR = `hc;
                12'd553: toneR = `hc;
                12'd554: toneR = `hc;
                12'd555: toneR = `hc;
                12'd556: toneR = `hc;
                12'd557: toneR = `hc;
                12'd558: toneR = `hc;
                12'd559: toneR = `hc;
                12'd560: toneR = `b;
                12'd561: toneR = `b;
                12'd562: toneR = `b;
                12'd563: toneR = `b;
                12'd564: toneR = `b;
                12'd565: toneR = `b;
                12'd566: toneR = `b;
                12'd567: toneR = `b;
                12'd568: toneR = `a;
                12'd569: toneR = `a;
                12'd570: toneR = `a;
                12'd571: toneR = `a;
                12'd572: toneR = `a;
                12'd573: toneR = `a;
                12'd574: toneR = `a;
                12'd575: toneR = `a;
                12'd576: toneR = `g;
                12'd577: toneR = `g;
                12'd578: toneR = `g;
                12'd579: toneR = `g;
                12'd580: toneR = `g;
                12'd581: toneR = `g;
                12'd582: toneR = `g;
                12'd583: toneR = `g;
                12'd584: toneR = `g;
                12'd585: toneR = `g;
                12'd586: toneR = `g;
                12'd587: toneR = `g;
                12'd588: toneR = `g;
                12'd589: toneR = `g;
                12'd590: toneR = `g;
                12'd591: toneR = `g;
                12'd592: toneR = `f;
                12'd593: toneR = `f;
                12'd594: toneR = `f;
                12'd595: toneR = `f;
                12'd596: toneR = `f;
                12'd597: toneR = `f;
                12'd598: toneR = `f;
                12'd599: toneR = `f;
                12'd600: toneR = `f;
                12'd601: toneR = `f;
                12'd602: toneR = `f;
                12'd603: toneR = `f;
                12'd604: toneR = `f;
                12'd605: toneR = `f;
                12'd606: toneR = `f;
                12'd607: toneR = `f;
                12'd608: toneR = `sil;
                12'd609: toneR = `sil;
                12'd610: toneR = `sil;
                12'd611: toneR = `sil;
                12'd612: toneR = `sil;
                12'd613: toneR = `sil;
                12'd614: toneR = `sil;
                12'd615: toneR = `sil;
                12'd616: toneR = `sil;
                12'd617: toneR = `sil;
                12'd618: toneR = `sil;
                12'd619: toneR = `sil;
                12'd620: toneR = `sil;
                12'd621: toneR = `sil;
                12'd622: toneR = `sil;
                12'd623: toneR = `sil;
                12'd624: toneR = `d;
                12'd625: toneR = `d;
                12'd626: toneR = `d;
                12'd627: toneR = `d;
                12'd628: toneR = `d;
                12'd629: toneR = `d;
                12'd630: toneR = `d;
                12'd631: toneR = `sil;
                12'd632: toneR = `d;
                12'd633: toneR = `d;
                12'd634: toneR = `d;
                12'd635: toneR = `d;
                12'd636: toneR = `d;
                12'd637: toneR = `d;
                12'd638: toneR = `d;
                12'd639: toneR = `d;
                12'd640: toneR = `e;
                12'd641: toneR = `e;
                12'd642: toneR = `e;
                12'd643: toneR = `e;
                12'd644: toneR = `e;
                12'd645: toneR = `e;
                12'd646: toneR = `e;
                12'd647: toneR = `e;
                12'd648: toneR = `f;
                12'd649: toneR = `f;
                12'd650: toneR = `f;
                12'd651: toneR = `f;
                12'd652: toneR = `f;
                12'd653: toneR = `f;
                12'd654: toneR = `f;
                12'd655: toneR = `f;
                12'd656: toneR = `lb;
                12'd657: toneR = `lb;
                12'd658: toneR = `lb;
                12'd659: toneR = `lb;
                12'd660: toneR = `lb;
                12'd661: toneR = `lb;
                12'd662: toneR = `lb;
                12'd663: toneR = `lb;
                12'd664: toneR = `b;
                12'd665: toneR = `b;
                12'd666: toneR = `b;
                12'd667: toneR = `b;
                12'd668: toneR = `b;
                12'd669: toneR = `b;
                12'd670: toneR = `b;
                12'd671: toneR = `b;
                12'd672: toneR = `a;
                12'd673: toneR = `a;
                12'd674: toneR = `a;
                12'd675: toneR = `a;
                12'd676: toneR = `a;
                12'd677: toneR = `a;
                12'd678: toneR = `a;
                12'd679: toneR = `a;
                12'd680: toneR = `g;
                12'd681: toneR = `g;
                12'd682: toneR = `g;
                12'd683: toneR = `g;
                12'd684: toneR = `g;
                12'd685: toneR = `g;
                12'd686: toneR = `g;
                12'd687: toneR = `g;
                12'd688: toneR = `a;
                12'd689: toneR = `a;
                12'd690: toneR = `a;
                12'd691: toneR = `a;
                12'd692: toneR = `a;
                12'd693: toneR = `a;
                12'd694: toneR = `a;
                12'd695: toneR = `a;
                12'd696: toneR = `a;
                12'd697: toneR = `a;
                12'd698: toneR = `a;
                12'd699: toneR = `a;
                12'd700: toneR = `a;
                12'd701: toneR = `a;
                12'd702: toneR = `a;
                12'd703: toneR = `a;
                12'd704: toneR = `g;
                12'd705: toneR = `g;
                12'd706: toneR = `g;
                12'd707: toneR = `g;
                12'd708: toneR = `g;
                12'd709: toneR = `g;
                12'd710: toneR = `g;
                12'd711: toneR = `g;
                12'd712: toneR = `g;
                12'd713: toneR = `g;
                12'd714: toneR = `g;
                12'd715: toneR = `g;
                12'd716: toneR = `g;
                12'd717: toneR = `g;
                12'd718: toneR = `g;
                12'd719: toneR = `g;
                12'd720: toneR = `sil;
                12'd721: toneR = `sil;
                12'd722: toneR = `sil;
                12'd723: toneR = `sil;
                12'd724: toneR = `sil;
                12'd725: toneR = `sil;
                12'd726: toneR = `sil;
                12'd727: toneR = `sil;
                12'd728: toneR = `sil;
                12'd729: toneR = `sil;
                12'd730: toneR = `sil;
                12'd731: toneR = `sil;
                12'd732: toneR = `sil;
                12'd733: toneR = `sil;
                12'd734: toneR = `sil;
                12'd735: toneR = `sil;
                12'd736: toneR = `e;
                12'd737: toneR = `e;
                12'd738: toneR = `e;
                12'd739: toneR = `e;
                12'd740: toneR = `e;
                12'd741: toneR = `e;
                12'd742: toneR = `e;
                12'd743: toneR = `sil;
                12'd744: toneR = `e;
                12'd745: toneR = `e;
                12'd746: toneR = `e;
                12'd747: toneR = `e;
                12'd748: toneR = `e;
                12'd749: toneR = `e;
                12'd750: toneR = `e;
                12'd751: toneR = `e;
                12'd752: toneR = `f;
                12'd753: toneR = `f;
                12'd754: toneR = `f;
                12'd755: toneR = `f;
                12'd756: toneR = `f;
                12'd757: toneR = `f;
                12'd758: toneR = `f;
                12'd759: toneR = `f;
                12'd760: toneR = `g;
                12'd761: toneR = `g;
                12'd762: toneR = `g;
                12'd763: toneR = `g;
                12'd764: toneR = `g;
                12'd765: toneR = `g;
                12'd766: toneR = `g;
                12'd767: toneR = `g;
                12'd768: toneR = `c;
                12'd769: toneR = `c;
                12'd770: toneR = `c;
                12'd771: toneR = `c;
                12'd772: toneR = `c;
                12'd773: toneR = `c;
                12'd774: toneR = `c;
                12'd775: toneR = `c;
                12'd776: toneR = `hc;
                12'd777: toneR = `hc;
                12'd778: toneR = `hc;
                12'd779: toneR = `hc;
                12'd780: toneR = `hc;
                12'd781: toneR = `hc;
                12'd782: toneR = `hc;
                12'd783: toneR = `hc;
                12'd784: toneR = `b;
                12'd785: toneR = `b;
                12'd786: toneR = `b;
                12'd787: toneR = `b;
                12'd788: toneR = `b;
                12'd789: toneR = `b;
                12'd790: toneR = `b;
                12'd791: toneR = `b;
                12'd792: toneR = `a;
                12'd793: toneR = `a;
                12'd794: toneR = `a;
                12'd795: toneR = `a;
                12'd796: toneR = `a;
                12'd797: toneR = `a;
                12'd798: toneR = `a;
                12'd799: toneR = `a;
                12'd800: toneR = `g;
                12'd801: toneR = `g;
                12'd802: toneR = `g;
                12'd803: toneR = `g;
                12'd804: toneR = `g;
                12'd805: toneR = `g;
                12'd806: toneR = `g;
                12'd807: toneR = `g;
                12'd808: toneR = `g;
                12'd809: toneR = `g;
                12'd810: toneR = `g;
                12'd811: toneR = `g;
                12'd812: toneR = `g;
                12'd813: toneR = `g;
                12'd814: toneR = `g;
                12'd815: toneR = `g;
                12'd816: toneR = `f;
                12'd817: toneR = `f;
                12'd818: toneR = `f;
                12'd819: toneR = `f;
                12'd820: toneR = `f;
                12'd821: toneR = `f;
                12'd822: toneR = `f;
                12'd823: toneR = `f;
                12'd824: toneR = `f;
                12'd825: toneR = `f;
                12'd826: toneR = `f;
                12'd827: toneR = `f;
                12'd828: toneR = `f;
                12'd829: toneR = `f;
                12'd830: toneR = `f;
                12'd831: toneR = `sil;
                12'd832: toneR = `f;
                12'd833: toneR = `f;
                12'd834: toneR = `f;
                12'd835: toneR = `f;
                12'd836: toneR = `f;
                12'd837: toneR = `f;
                12'd838: toneR = `f;
                12'd839: toneR = `f;
                12'd840: toneR = `g;
                12'd841: toneR = `g;
                12'd842: toneR = `g;
                12'd843: toneR = `g;
                12'd844: toneR = `g;
                12'd845: toneR = `g;
                12'd846: toneR = `g;
                12'd847: toneR = `g;
                12'd848: toneR = `a;
                12'd849: toneR = `a;
                12'd850: toneR = `a;
                12'd851: toneR = `a;
                12'd852: toneR = `a;
                12'd853: toneR = `a;
                12'd854: toneR = `a;
                12'd855: toneR = `a;
                12'd856: toneR = `b;
                12'd857: toneR = `b;
                12'd858: toneR = `b;
                12'd859: toneR = `b;
                12'd860: toneR = `b;
                12'd861: toneR = `b;
                12'd862: toneR = `b;
                12'd863: toneR = `b;
                12'd864: toneR = `sil;
                12'd865: toneR = `sil;
                12'd866: toneR = `sil;
                12'd867: toneR = `sil;
                12'd868: toneR = `sil;
                12'd869: toneR = `sil;
                12'd870: toneR = `sil;
                12'd871: toneR = `sil;
                12'd872: toneR = `g;
                12'd873: toneR = `g;
                12'd874: toneR = `g;
                12'd875: toneR = `g;
                12'd876: toneR = `g;
                12'd877: toneR = `g;
                12'd878: toneR = `g;
                12'd879: toneR = `g;
                12'd880: toneR = `g;
                12'd881: toneR = `g;
                12'd882: toneR = `g;
                12'd883: toneR = `g;
                12'd884: toneR = `g;
                12'd885: toneR = `g;
                12'd886: toneR = `g;
                12'd887: toneR = `g;
                12'd888: toneR = `a;
                12'd889: toneR = `a;
                12'd890: toneR = `a;
                12'd891: toneR = `a;
                12'd892: toneR = `a;
                12'd893: toneR = `a;
                12'd894: toneR = `a;
                12'd895: toneR = `a;
                12'd896: toneR = `a;
                12'd897: toneR = `a;
                12'd898: toneR = `a;
                12'd899: toneR = `a;
                12'd900: toneR = `a;
                12'd901: toneR = `a;
                12'd902: toneR = `a;
                12'd903: toneR = `a;
                12'd904: toneR = `b;
                12'd905: toneR = `b;
                12'd906: toneR = `b;
                12'd907: toneR = `b;
                12'd908: toneR = `b;
                12'd909: toneR = `b;
                12'd910: toneR = `b;
                12'd911: toneR = `b;
                12'd912: toneR = `b;
                12'd913: toneR = `b;
                12'd914: toneR = `b;
                12'd915: toneR = `b;
                12'd916: toneR = `b;
                12'd917: toneR = `b;
                12'd918: toneR = `b;
                12'd919: toneR = `b;
                12'd920: toneR = `hc;
                12'd921: toneR = `hc;
                12'd922: toneR = `hc;
                12'd923: toneR = `hc;
                12'd924: toneR = `hc;
                12'd925: toneR = `hc;
                12'd926: toneR = `hc;
                12'd927: toneR = `hc;
                12'd928: toneR = `hc;
                12'd929: toneR = `hc;
                12'd930: toneR = `hc;
                12'd931: toneR = `hc;
                12'd932: toneR = `hc;
                12'd933: toneR = `hc;
                12'd934: toneR = `hc;
                12'd935: toneR = `hc;
                12'd936: toneR = `hc;
                12'd937: toneR = `hc;
                12'd938: toneR = `hc;
                12'd939: toneR = `hc;
                12'd940: toneR = `hc;
                12'd941: toneR = `hc;
                12'd942: toneR = `hc;
                12'd943: toneR = `hc;
                12'd944: toneR = `hc;
                12'd945: toneR = `hc;
                12'd946: toneR = `hc;
                12'd947: toneR = `hc;
                12'd948: toneR = `hc;
                12'd949: toneR = `hc;
                12'd950: toneR = `hc;
                12'd951: toneR = `hc;
                12'd952: toneR = `hc;
                12'd953: toneR = `hc;
                12'd954: toneR = `hc;
                12'd955: toneR = `hc;
                12'd956: toneR = `hc;
                12'd957: toneR = `hc;
                12'd958: toneR = `hc;
                12'd959: toneR = `hc;
                12'd960: toneR = `sil;
                12'd961: toneR = `sil;
                12'd962: toneR = `sil;
                12'd963: toneR = `sil;
                12'd964: toneR = `sil;
                12'd965: toneR = `sil;
                12'd966: toneR = `sil;
                12'd967: toneR = `sil;
                12'd968: toneR = `sil;
                12'd969: toneR = `sil;
                12'd970: toneR = `sil;
                12'd971: toneR = `sil;
                12'd972: toneR = `sil;
                12'd973: toneR = `sil;
                12'd974: toneR = `sil;
                12'd975: toneR = `sil;
                12'd976: toneR = `sil;
                12'd977: toneR = `sil;
                12'd978: toneR = `sil;
                12'd979: toneR = `sil;
                12'd980: toneR = `sil;
                12'd981: toneR = `sil;
                12'd982: toneR = `sil;
                12'd983: toneR = `sil;
                12'd984: toneR = `hc;
                12'd985: toneR = `hc;
                12'd986: toneR = `hc;
                12'd987: toneR = `hc;
                12'd988: toneR = `hc;
                12'd989: toneR = `hc;
                12'd990: toneR = `hc;
                12'd991: toneR = `hc;
                12'd992: toneR = `b;
                12'd993: toneR = `b;
                12'd994: toneR = `b;
                12'd995: toneR = `b;
                12'd996: toneR = `b;
                12'd997: toneR = `b;
                12'd998: toneR = `b;
                12'd999: toneR = `b;
                12'd1000: toneR = `sa;
                12'd1001: toneR = `sa;
                12'd1002: toneR = `sa;
                12'd1003: toneR = `sa;
                12'd1004: toneR = `sa;
                12'd1005: toneR = `sa;
                12'd1006: toneR = `sa;
                12'd1007: toneR = `sa;
                12'd1008: toneR = `a;
                12'd1009: toneR = `a;
                12'd1010: toneR = `a;
                12'd1011: toneR = `a;
                12'd1012: toneR = `a;
                12'd1013: toneR = `a;
                12'd1014: toneR = `a;
                12'd1015: toneR = `a;
                12'd1016: toneR = `a;
                12'd1017: toneR = `a;
                12'd1018: toneR = `a;
                12'd1019: toneR = `a;
                12'd1020: toneR = `a;
                12'd1021: toneR = `a;
                12'd1022: toneR = `a;
                12'd1023: toneR = `a;
                12'd1024: toneR = `hc;
                12'd1025: toneR = `hc;
                12'd1026: toneR = `hc;
                12'd1027: toneR = `hc;
                12'd1028: toneR = `hc;
                12'd1029: toneR = `hc;
                12'd1030: toneR = `hc;
                12'd1031: toneR = `hc;
                12'd1032: toneR = `hc;
                12'd1033: toneR = `hc;
                12'd1034: toneR = `hc;
                12'd1035: toneR = `hc;
                12'd1036: toneR = `hc;
                12'd1037: toneR = `hc;
                12'd1038: toneR = `hc;
                12'd1039: toneR = `hc;
                12'd1040: toneR = `hd;
                12'd1041: toneR = `hd;
                12'd1042: toneR = `hd;
                12'd1043: toneR = `hd;
                12'd1044: toneR = `hd;
                12'd1045: toneR = `hd;
                12'd1046: toneR = `hd;
                12'd1047: toneR = `hd;
                12'd1048: toneR = `hd;
                12'd1049: toneR = `hd;
                12'd1050: toneR = `hd;
                12'd1051: toneR = `hd;
                12'd1052: toneR = `hd;
                12'd1053: toneR = `hd;
                12'd1054: toneR = `hd;
                12'd1055: toneR = `hd;
                12'd1056: toneR = `hc;
                12'd1057: toneR = `hc;
                12'd1058: toneR = `hc;
                12'd1059: toneR = `hc;
                12'd1060: toneR = `hc;
                12'd1061: toneR = `hc;
                12'd1062: toneR = `hc;
                12'd1063: toneR = `hc;
                12'd1064: toneR = `hc;
                12'd1065: toneR = `hc;
                12'd1066: toneR = `hc;
                12'd1067: toneR = `hc;
                12'd1068: toneR = `hc;
                12'd1069: toneR = `hc;
                12'd1070: toneR = `hc;
                12'd1071: toneR = `hc;
                12'd1072: toneR = `g;
                12'd1073: toneR = `g;
                12'd1074: toneR = `g;
                12'd1075: toneR = `g;
                12'd1076: toneR = `g;
                12'd1077: toneR = `g;
                12'd1078: toneR = `g;
                12'd1079: toneR = `g;
                12'd1080: toneR = `g;
                12'd1081: toneR = `g;
                12'd1082: toneR = `g;
                12'd1083: toneR = `g;
                12'd1084: toneR = `g;
                12'd1085: toneR = `g;
                12'd1086: toneR = `g;
                12'd1087: toneR = `g;
                12'd1088: toneR = `sil;
                12'd1089: toneR = `sil;
                12'd1090: toneR = `sil;
                12'd1091: toneR = `sil;
                12'd1092: toneR = `sil;
                12'd1093: toneR = `sil;
                12'd1094: toneR = `sil;
                12'd1095: toneR = `sil;
                12'd1096: toneR = `sil;
                12'd1097: toneR = `sil;
                12'd1098: toneR = `sil;
                12'd1099: toneR = `sil;
                12'd1100: toneR = `sil;
                12'd1101: toneR = `sil;
                12'd1102: toneR = `sil;
                12'd1103: toneR = `sil;
                12'd1104: toneR = `sil;
                12'd1105: toneR = `sil;
                12'd1106: toneR = `sil;
                12'd1107: toneR = `sil;
                12'd1108: toneR = `sil;
                12'd1109: toneR = `sil;
                12'd1110: toneR = `sil;
                12'd1111: toneR = `sil;
                12'd1112: toneR = `hc;
                12'd1113: toneR = `hc;
                12'd1114: toneR = `hc;
                12'd1115: toneR = `hc;
                12'd1116: toneR = `hc;
                12'd1117: toneR = `hc;
                12'd1118: toneR = `hc;
                12'd1119: toneR = `hc;
                12'd1120: toneR = `b;
                12'd1121: toneR = `b;
                12'd1122: toneR = `b;
                12'd1123: toneR = `b;
                12'd1124: toneR = `b;
                12'd1125: toneR = `b;
                12'd1126: toneR = `b;
                12'd1127: toneR = `b;
                12'd1128: toneR = `sa;
                12'd1129: toneR = `sa;
                12'd1130: toneR = `sa;
                12'd1131: toneR = `sa;
                12'd1132: toneR = `sa;
                12'd1133: toneR = `sa;
                12'd1134: toneR = `sa;
                12'd1135: toneR = `sa;
                12'd1136: toneR = `a;
                12'd1137: toneR = `a;
                12'd1138: toneR = `a;
                12'd1139: toneR = `a;
                12'd1140: toneR = `a;
                12'd1141: toneR = `a;
                12'd1142: toneR = `a;
                12'd1143: toneR = `a;
                12'd1144: toneR = `a;
                12'd1145: toneR = `a;
                12'd1146: toneR = `a;
                12'd1147: toneR = `a;
                12'd1148: toneR = `a;
                12'd1149: toneR = `a;
                12'd1150: toneR = `a;
                12'd1151: toneR = `a;
                12'd1152: toneR = `hc;
                12'd1153: toneR = `hc;
                12'd1154: toneR = `hc;
                12'd1155: toneR = `hc;
                12'd1156: toneR = `hc;
                12'd1157: toneR = `hc;
                12'd1158: toneR = `hc;
                12'd1159: toneR = `hc;
                12'd1160: toneR = `hc;
                12'd1161: toneR = `hc;
                12'd1162: toneR = `hc;
                12'd1163: toneR = `hc;
                12'd1164: toneR = `hc;
                12'd1165: toneR = `hc;
                12'd1166: toneR = `hc;
                12'd1167: toneR = `hc;
                12'd1168: toneR = `hd;
                12'd1169: toneR = `hd;
                12'd1170: toneR = `hd;
                12'd1171: toneR = `hd;
                12'd1172: toneR = `hd;
                12'd1173: toneR = `hd;
                12'd1174: toneR = `hd;
                12'd1175: toneR = `hd;
                12'd1176: toneR = `hd;
                12'd1177: toneR = `hd;
                12'd1178: toneR = `hd;
                12'd1179: toneR = `hd;
                12'd1180: toneR = `hd;
                12'd1181: toneR = `hd;
                12'd1182: toneR = `hd;
                12'd1183: toneR = `hd;
                12'd1184: toneR = `hc;
                12'd1185: toneR = `hc;
                12'd1186: toneR = `hc;
                12'd1187: toneR = `hc;
                12'd1188: toneR = `hc;
                12'd1189: toneR = `hc;
                12'd1190: toneR = `hc;
                12'd1191: toneR = `hc;
                12'd1192: toneR = `hc;
                12'd1193: toneR = `hc;
                12'd1194: toneR = `hc;
                12'd1195: toneR = `hc;
                12'd1196: toneR = `hc;
                12'd1197: toneR = `hc;
                12'd1198: toneR = `hc;
                12'd1199: toneR = `hc;
                12'd1200: toneR = `g;
                12'd1201: toneR = `g;
                12'd1202: toneR = `g;
                12'd1203: toneR = `g;
                12'd1204: toneR = `g;
                12'd1205: toneR = `g;
                12'd1206: toneR = `g;
                12'd1207: toneR = `g;
                12'd1208: toneR = `g;
                12'd1209: toneR = `g;
                12'd1210: toneR = `g;
                12'd1211: toneR = `g;
                12'd1212: toneR = `g;
                12'd1213: toneR = `g;
                12'd1214: toneR = `g;
                12'd1215: toneR = `g;
                12'd1216: toneR = `sil;
                12'd1217: toneR = `sil;
                12'd1218: toneR = `sil;
                12'd1219: toneR = `sil;
                12'd1220: toneR = `sil;
                12'd1221: toneR = `sil;
                12'd1222: toneR = `sil;
                12'd1223: toneR = `sil;
                12'd1224: toneR = `sil;
                12'd1225: toneR = `sil;
                12'd1226: toneR = `sil;
                12'd1227: toneR = `sil;
                12'd1228: toneR = `sil;
                12'd1229: toneR = `sil;
                12'd1230: toneR = `sil;
                12'd1231: toneR = `sil;
                12'd1232: toneR = `sil;
                12'd1233: toneR = `sil;
                12'd1234: toneR = `sil;
                12'd1235: toneR = `sil;
                12'd1236: toneR = `sil;
                12'd1237: toneR = `sil;
                12'd1238: toneR = `sil;
                12'd1239: toneR = `sil;
                12'd1240: toneR = `hc;
                12'd1241: toneR = `hc;
                12'd1242: toneR = `hc;
                12'd1243: toneR = `hc;
                12'd1244: toneR = `hc;
                12'd1245: toneR = `hc;
                12'd1246: toneR = `hc;
                12'd1247: toneR = `hc;
                12'd1248: toneR = `b;
                12'd1249: toneR = `b;
                12'd1250: toneR = `b;
                12'd1251: toneR = `b;
                12'd1252: toneR = `b;
                12'd1253: toneR = `b;
                12'd1254: toneR = `b;
                12'd1255: toneR = `b;
                12'd1256: toneR = `sa;
                12'd1257: toneR = `sa;
                12'd1258: toneR = `sa;
                12'd1259: toneR = `sa;
                12'd1260: toneR = `sa;
                12'd1261: toneR = `sa;
                12'd1262: toneR = `sa;
                12'd1263: toneR = `sa;
                12'd1264: toneR = `a;
                12'd1265: toneR = `a;
                12'd1266: toneR = `a;
                12'd1267: toneR = `a;
                12'd1268: toneR = `a;
                12'd1269: toneR = `a;
                12'd1270: toneR = `a;
                12'd1271: toneR = `a;
                12'd1272: toneR = `a;
                12'd1273: toneR = `a;
                12'd1274: toneR = `a;
                12'd1275: toneR = `a;
                12'd1276: toneR = `a;
                12'd1277: toneR = `a;
                12'd1278: toneR = `a;
                12'd1279: toneR = `a;
                12'd1280: toneR = `hc;
                12'd1281: toneR = `hc;
                12'd1282: toneR = `hc;
                12'd1283: toneR = `hc;
                12'd1284: toneR = `hc;
                12'd1285: toneR = `hc;
                12'd1286: toneR = `hc;
                12'd1287: toneR = `hc;
                12'd1288: toneR = `hc;
                12'd1289: toneR = `hc;
                12'd1290: toneR = `hc;
                12'd1291: toneR = `hc;
                12'd1292: toneR = `hc;
                12'd1293: toneR = `hc;
                12'd1294: toneR = `hc;
                12'd1295: toneR = `hc;
                12'd1296: toneR = `hd;
                12'd1297: toneR = `hd;
                12'd1298: toneR = `hd;
                12'd1299: toneR = `hd;
                12'd1300: toneR = `hd;
                12'd1301: toneR = `hd;
                12'd1302: toneR = `hd;
                12'd1303: toneR = `hd;
                12'd1304: toneR = `hd;
                12'd1305: toneR = `hd;
                12'd1306: toneR = `hd;
                12'd1307: toneR = `hd;
                12'd1308: toneR = `hd;
                12'd1309: toneR = `hd;
                12'd1310: toneR = `hd;
                12'd1311: toneR = `hd;
                12'd1312: toneR = `hc;
                12'd1313: toneR = `hc;
                12'd1314: toneR = `hc;
                12'd1315: toneR = `hc;
                12'd1316: toneR = `hc;
                12'd1317: toneR = `hc;
                12'd1318: toneR = `hc;
                12'd1319: toneR = `hc;
                12'd1320: toneR = `hd;
                12'd1321: toneR = `hd;
                12'd1322: toneR = `hd;
                12'd1323: toneR = `hd;
                12'd1324: toneR = `hd;
                12'd1325: toneR = `hd;
                12'd1326: toneR = `hd;
                12'd1327: toneR = `hd;
                12'd1328: toneR = `he;
                12'd1329: toneR = `he;
                12'd1330: toneR = `he;
                12'd1331: toneR = `he;
                12'd1332: toneR = `he;
                12'd1333: toneR = `he;
                12'd1334: toneR = `he;
                12'd1335: toneR = `he;
                12'd1336: toneR = `hd;
                12'd1337: toneR = `hd;
                12'd1338: toneR = `hd;
                12'd1339: toneR = `hd;
                12'd1340: toneR = `hd;
                12'd1341: toneR = `hd;
                12'd1342: toneR = `hd;
                12'd1343: toneR = `hd;
                12'd1344: toneR = `he;
                12'd1345: toneR = `he;
                12'd1346: toneR = `he;
                12'd1347: toneR = `he;
                12'd1348: toneR = `he;
                12'd1349: toneR = `he;
                12'd1350: toneR = `he;
                12'd1351: toneR = `he;
                12'd1352: toneR = `hc;
                12'd1353: toneR = `hc;
                12'd1354: toneR = `hc;
                12'd1355: toneR = `hc;
                12'd1356: toneR = `hc;
                12'd1357: toneR = `hc;
                12'd1358: toneR = `hc;
                12'd1359: toneR = `hc;
                12'd1360: toneR = `sil;
                12'd1361: toneR = `sil;
                12'd1362: toneR = `sil;
                12'd1363: toneR = `sil;
                12'd1364: toneR = `sil;
                12'd1365: toneR = `sil;
                12'd1366: toneR = `sil;
                12'd1367: toneR = `sil;
                12'd1368: toneR = `hc;
                12'd1369: toneR = `hc;
                12'd1370: toneR = `hc;
                12'd1371: toneR = `hc;
                12'd1372: toneR = `hc;
                12'd1373: toneR = `hc;
                12'd1374: toneR = `hc;
                12'd1375: toneR = `hc;
                12'd1376: toneR = `hd;
                12'd1377: toneR = `hd;
                12'd1378: toneR = `hd;
                12'd1379: toneR = `hd;
                12'd1380: toneR = `hd;
                12'd1381: toneR = `hd;
                12'd1382: toneR = `hd;
                12'd1383: toneR = `hd;
                12'd1384: toneR = `he;
                12'd1385: toneR = `he;
                12'd1386: toneR = `he;
                12'd1387: toneR = `he;
                12'd1388: toneR = `he;
                12'd1389: toneR = `he;
                12'd1390: toneR = `he;
                12'd1391: toneR = `he;
                12'd1392: toneR = `hf;
                12'd1393: toneR = `hf;
                12'd1394: toneR = `hf;
                12'd1395: toneR = `hf;
                12'd1396: toneR = `hf;
                12'd1397: toneR = `hf;
                12'd1398: toneR = `hf;
                12'd1399: toneR = `hf;
                12'd1400: toneR = `hf;
                12'd1401: toneR = `hf;
                12'd1402: toneR = `hf;
                12'd1403: toneR = `hf;
                12'd1404: toneR = `hf;
                12'd1405: toneR = `hf;
                12'd1406: toneR = `hf;
                12'd1407: toneR = `hf;
                12'd1408: toneR = `a;
                12'd1409: toneR = `a;
                12'd1410: toneR = `a;
                12'd1411: toneR = `a;
                12'd1412: toneR = `a;
                12'd1413: toneR = `a;
                12'd1414: toneR = `a;
                12'd1415: toneR = `a;
                12'd1416: toneR = `a;
                12'd1417: toneR = `a;
                12'd1418: toneR = `a;
                12'd1419: toneR = `a;
                12'd1420: toneR = `a;
                12'd1421: toneR = `a;
                12'd1422: toneR = `a;
                12'd1423: toneR = `a;
                12'd1424: toneR = `b;
                12'd1425: toneR = `b;
                12'd1426: toneR = `b;
                12'd1427: toneR = `b;
                12'd1428: toneR = `b;
                12'd1429: toneR = `b;
                12'd1430: toneR = `b;
                12'd1431: toneR = `b;
                12'd1432: toneR = `b;
                12'd1433: toneR = `b;
                12'd1434: toneR = `b;
                12'd1435: toneR = `b;
                12'd1436: toneR = `b;
                12'd1437: toneR = `b;
                12'd1438: toneR = `b;
                12'd1439: toneR = `b;
                12'd1440: toneR = `hd;
                12'd1441: toneR = `hd;
                12'd1442: toneR = `hd;
                12'd1443: toneR = `hd;
                12'd1444: toneR = `hd;
                12'd1445: toneR = `hd;
                12'd1446: toneR = `hd;
                12'd1447: toneR = `hd;
                12'd1448: toneR = `hd;
                12'd1449: toneR = `hd;
                12'd1450: toneR = `hd;
                12'd1451: toneR = `hd;
                12'd1452: toneR = `hd;
                12'd1453: toneR = `hd;
                12'd1454: toneR = `hd;
                12'd1455: toneR = `hd;
                12'd1456: toneR = `hc;
                12'd1457: toneR = `hc;
                12'd1458: toneR = `hc;
                12'd1459: toneR = `hc;
                12'd1460: toneR = `hc;
                12'd1461: toneR = `hc;
                12'd1462: toneR = `hc;
                12'd1463: toneR = `hc;
                12'd1464: toneR = `hc;
                12'd1465: toneR = `hc;
                12'd1466: toneR = `hc;
                12'd1467: toneR = `hc;
                12'd1468: toneR = `hc;
                12'd1469: toneR = `hc;
                12'd1470: toneR = `hc;
                12'd1471: toneR = `hc;
                12'd1472: toneR = `sil;
                12'd1473: toneR = `sil;
                12'd1474: toneR = `sil;
                12'd1475: toneR = `sil;
                12'd1476: toneR = `sil;
                12'd1477: toneR = `sil;
                12'd1478: toneR = `sil;
                12'd1479: toneR = `sil;
                12'd1480: toneR = `sil;
                12'd1481: toneR = `sil;
                12'd1482: toneR = `sil;
                12'd1483: toneR = `sil;
                12'd1484: toneR = `sil;
                12'd1485: toneR = `sil;
                12'd1486: toneR = `sil;
                12'd1487: toneR = `sil;
                12'd1488: toneR = `sil;
                12'd1489: toneR = `sil;
                12'd1490: toneR = `sil;
                12'd1491: toneR = `sil;
                12'd1492: toneR = `sil;
                12'd1493: toneR = `sil;
                12'd1494: toneR = `sil;
                12'd1495: toneR = `sil;
                12'd1496: toneR = `sil;
                12'd1497: toneR = `sil;
                12'd1498: toneR = `sil;
                12'd1499: toneR = `sil;
                12'd1500: toneR = `sil;
                12'd1501: toneR = `sil;
                12'd1502: toneR = `sil;
                12'd1503: toneR = `sil;
                12'd1504: toneR = `sil;
                12'd1505: toneR = `sil;
                12'd1506: toneR = `sil;
                12'd1507: toneR = `sil;
                12'd1508: toneR = `sil;
                12'd1509: toneR = `sil;
                12'd1510: toneR = `sil;
                12'd1511: toneR = `sil;
                12'd1512: toneR = `sil;
                12'd1513: toneR = `sil;
                12'd1514: toneR = `sil;
                12'd1515: toneR = `sil;
                12'd1516: toneR = `sil;
                12'd1517: toneR = `sil;
                12'd1518: toneR = `sil;
                12'd1519: toneR = `sil;
                12'd1520: toneR = `sil;
                12'd1521: toneR = `sil;
                12'd1522: toneR = `sil;
                12'd1523: toneR = `sil;
                12'd1524: toneR = `sil;
                12'd1525: toneR = `sil;
                12'd1526: toneR = `sil;
                12'd1527: toneR = `sil;
                12'd1528: toneR = `sil;
                12'd1529: toneR = `sil;
                12'd1530: toneR = `sil;
                12'd1531: toneR = `sil;
                12'd1532: toneR = `sil;
                12'd1533: toneR = `sil;
                12'd1534: toneR = `sil;
                12'd1535: toneR = `sil;
            default:toneR = `sil;
        endcase
    end
    else toneR = `sil;
end

always @(*) begin
    if(en) begin
        case(ibeatNum)
                12'd0: toneL = `sil;
                12'd1: toneL = `sil;
                12'd2: toneL = `sil;
                12'd3: toneL = `sil;
                12'd4: toneL = `sil;
                12'd5: toneL = `sil;
                12'd6: toneL = `sil;
                12'd7: toneL = `sil;
                12'd8: toneL = `sil;
                12'd9: toneL = `sil;
                12'd10: toneL = `sil;
                12'd11: toneL = `sil;
                12'd12: toneL = `sil;
                12'd13: toneL = `sil;
                12'd14: toneL = `sil;
                12'd15: toneL = `sil;
                12'd16: toneL = `sil;
                12'd17: toneL = `sil;
                12'd18: toneL = `sil;
                12'd19: toneL = `sil;
                12'd20: toneL = `sil;
                12'd21: toneL = `sil;
                12'd22: toneL = `sil;
                12'd23: toneL = `sil;
                12'd24: toneL = `lg;
                12'd25: toneL = `lg;
                12'd26: toneL = `lg;
                12'd27: toneL = `lg;
                12'd28: toneL = `sil;
                12'd29: toneL = `sil;
                12'd30: toneL = `sil;
                12'd31: toneL = `sil;
                12'd32: toneL = `sil;
                12'd33: toneL = `sil;
                12'd34: toneL = `sil;
                12'd35: toneL = `sil;
                12'd36: toneL = `sil;
                12'd37: toneL = `sil;
                12'd38: toneL = `sil;
                12'd39: toneL = `sil;
                12'd40: toneL = `sil;
                12'd41: toneL = `sil;
                12'd42: toneL = `sil;
                12'd43: toneL = `sil;
                12'd44: toneL = `sil;
                12'd45: toneL = `sil;
                12'd46: toneL = `sil;
                12'd47: toneL = `sil;
                12'd48: toneL = `sil;
                12'd49: toneL = `sil;
                12'd50: toneL = `sil;
                12'd51: toneL = `sil;
                12'd52: toneL = `sil;
                12'd53: toneL = `sil;
                12'd54: toneL = `sil;
                12'd55: toneL = `sil;
                12'd56: toneL = `lg;
                12'd57: toneL = `lg;
                12'd58: toneL = `lg;
                12'd59: toneL = `lg;
                12'd60: toneL = `sil;
                12'd61: toneL = `sil;
                12'd62: toneL = `sil;
                12'd63: toneL = `sil;
                12'd64: toneL = `d;
                12'd65: toneL = `d;
                12'd66: toneL = `d;
                12'd67: toneL = `d;
                12'd68: toneL = `d;
                12'd69: toneL = `d;
                12'd70: toneL = `d;
                12'd71: toneL = `d;
                12'd72: toneL = `d;
                12'd73: toneL = `d;
                12'd74: toneL = `d;
                12'd75: toneL = `d;
                12'd76: toneL = `d;
                12'd77: toneL = `d;
                12'd78: toneL = `d;
                12'd79: toneL = `d;
                12'd80: toneL = `e;
                12'd81: toneL = `e;
                12'd82: toneL = `e;
                12'd83: toneL = `e;
                12'd84: toneL = `e;
                12'd85: toneL = `e;
                12'd86: toneL = `e;
                12'd87: toneL = `e;
                12'd88: toneL = `e;
                12'd89: toneL = `e;
                12'd90: toneL = `e;
                12'd91: toneL = `e;
                12'd92: toneL = `e;
                12'd93: toneL = `e;
                12'd94: toneL = `e;
                12'd95: toneL = `e;
                12'd96: toneL = `f;
                12'd97: toneL = `f;
                12'd98: toneL = `f;
                12'd99: toneL = `f;
                12'd100: toneL = `f;
                12'd101: toneL = `f;
                12'd102: toneL = `f;
                12'd103: toneL = `f;
                12'd104: toneL = `f;
                12'd105: toneL = `f;
                12'd106: toneL = `f;
                12'd107: toneL = `f;
                12'd108: toneL = `f;
                12'd109: toneL = `f;
                12'd110: toneL = `f;
                12'd111: toneL = `f;
                12'd112: toneL = `g;
                12'd113: toneL = `g;
                12'd114: toneL = `g;
                12'd115: toneL = `g;
                12'd116: toneL = `g;
                12'd117: toneL = `g;
                12'd118: toneL = `g;
                12'd119: toneL = `g;
                12'd120: toneL = `g;
                12'd121: toneL = `g;
                12'd122: toneL = `g;
                12'd123: toneL = `g;
                12'd124: toneL = `g;
                12'd125: toneL = `g;
                12'd126: toneL = `g;
                12'd127: toneL = `g;
                12'd128: toneL = `g;
                12'd129: toneL = `g;
                12'd130: toneL = `g;
                12'd131: toneL = `g;
                12'd132: toneL = `g;
                12'd133: toneL = `g;
                12'd134: toneL = `g;
                12'd135: toneL = `g;
                12'd136: toneL = `g;
                12'd137: toneL = `g;
                12'd138: toneL = `g;
                12'd139: toneL = `g;
                12'd140: toneL = `g;
                12'd141: toneL = `g;
                12'd142: toneL = `g;
                12'd143: toneL = `sil;
                12'd144: toneL = `g;
                12'd145: toneL = `g;
                12'd146: toneL = `g;
                12'd147: toneL = `g;
                12'd148: toneL = `g;
                12'd149: toneL = `g;
                12'd150: toneL = `g;
                12'd151: toneL = `g;
                12'd152: toneL = `sf;
                12'd153: toneL = `sf;
                12'd154: toneL = `sf;
                12'd155: toneL = `sf;
                12'd156: toneL = `g;
                12'd157: toneL = `g;
                12'd158: toneL = `g;
                12'd159: toneL = `g;
                12'd160: toneL = `g;
                12'd161: toneL = `g;
                12'd162: toneL = `g;
                12'd163: toneL = `g;
                12'd164: toneL = `g;
                12'd165: toneL = `g;
                12'd166: toneL = `g;
                12'd167: toneL = `g;
                12'd168: toneL = `g;
                12'd169: toneL = `g;
                12'd170: toneL = `g;
                12'd171: toneL = `g;
                12'd172: toneL = `sil;
                12'd173: toneL = `sil;
                12'd174: toneL = `sil;
                12'd175: toneL = `sil;
                12'd176: toneL = `sil;
                12'd177: toneL = `sil;
                12'd178: toneL = `sil;
                12'd179: toneL = `sil;
                12'd180: toneL = `sil;
                12'd181: toneL = `sil;
                12'd182: toneL = `sil;
                12'd183: toneL = `sil;
                12'd184: toneL = `sil;
                12'd185: toneL = `sil;
                12'd186: toneL = `sil;
                12'd187: toneL = `sil;
                12'd188: toneL = `sil;
                12'd189: toneL = `sil;
                12'd190: toneL = `sil;
                12'd191: toneL = `sil;
                12'd192: toneL = `f;
                12'd193: toneL = `f;
                12'd194: toneL = `f;
                12'd195: toneL = `f;
                12'd196: toneL = `f;
                12'd197: toneL = `f;
                12'd198: toneL = `f;
                12'd199: toneL = `f;
                12'd200: toneL = `f;
                12'd201: toneL = `f;
                12'd202: toneL = `f;
                12'd203: toneL = `f;
                12'd204: toneL = `f;
                12'd205: toneL = `f;
                12'd206: toneL = `f;
                12'd207: toneL = `sil;
                12'd208: toneL = `f;
                12'd209: toneL = `f;
                12'd210: toneL = `f;
                12'd211: toneL = `f;
                12'd212: toneL = `f;
                12'd213: toneL = `f;
                12'd214: toneL = `f;
                12'd215: toneL = `f;
                12'd216: toneL = `g;
                12'd217: toneL = `g;
                12'd218: toneL = `g;
                12'd219: toneL = `g;
                12'd220: toneL = `d;
                12'd221: toneL = `d;
                12'd222: toneL = `d;
                12'd223: toneL = `d;
                12'd224: toneL = `d;
                12'd225: toneL = `d;
                12'd226: toneL = `d;
                12'd227: toneL = `d;
                12'd228: toneL = `d;
                12'd229: toneL = `d;
                12'd230: toneL = `d;
                12'd231: toneL = `d;
                12'd232: toneL = `d;
                12'd233: toneL = `d;
                12'd234: toneL = `d;
                12'd235: toneL = `d;
                12'd236: toneL = `sil;
                12'd237: toneL = `sil;
                12'd238: toneL = `sil;
                12'd239: toneL = `sil;
                12'd240: toneL = `la;
                12'd241: toneL = `la;
                12'd242: toneL = `la;
                12'd243: toneL = `la;
                12'd244: toneL = `la;
                12'd245: toneL = `la;
                12'd246: toneL = `la;
                12'd247: toneL = `la;
                12'd248: toneL = `lb;
                12'd249: toneL = `lb;
                12'd250: toneL = `lb;
                12'd251: toneL = `lb;
                12'd252: toneL = `lb;
                12'd253: toneL = `lb;
                12'd254: toneL = `lb;
                12'd255: toneL = `lb;
                12'd256: toneL = `c;
                12'd257: toneL = `c;
                12'd258: toneL = `c;
                12'd259: toneL = `c;
                12'd260: toneL = `c;
                12'd261: toneL = `c;
                12'd262: toneL = `c;
                12'd263: toneL = `c;
                12'd264: toneL = `c;
                12'd265: toneL = `c;
                12'd266: toneL = `c;
                12'd267: toneL = `c;
                12'd268: toneL = `c;
                12'd269: toneL = `c;
                12'd270: toneL = `c;
                12'd271: toneL = `c;
                12'd272: toneL = `c;
                12'd273: toneL = `c;
                12'd274: toneL = `c;
                12'd275: toneL = `c;
                12'd276: toneL = `c;
                12'd277: toneL = `c;
                12'd278: toneL = `c;
                12'd279: toneL = `c;
                12'd280: toneL = `c;
                12'd281: toneL = `c;
                12'd282: toneL = `c;
                12'd283: toneL = `c;
                12'd284: toneL = `c;
                12'd285: toneL = `c;
                12'd286: toneL = `c;
                12'd287: toneL = `c;
                12'd288: toneL = `sil;
                12'd289: toneL = `sil;
                12'd290: toneL = `sil;
                12'd291: toneL = `sil;
                12'd292: toneL = `sil;
                12'd293: toneL = `sil;
                12'd294: toneL = `sil;
                12'd295: toneL = `sil;
                12'd296: toneL = `sil;
                12'd297: toneL = `sil;
                12'd298: toneL = `sil;
                12'd299: toneL = `sil;
                12'd300: toneL = `sil;
                12'd301: toneL = `sil;
                12'd302: toneL = `sil;
                12'd303: toneL = `sil;
                12'd304: toneL = `sil;
                12'd305: toneL = `sil;
                12'd306: toneL = `sil;
                12'd307: toneL = `sil;
                12'd308: toneL = `sil;
                12'd309: toneL = `sil;
                12'd310: toneL = `sil;
                12'd311: toneL = `sil;
                12'd312: toneL = `lg;
                12'd313: toneL = `lg;
                12'd314: toneL = `lg;
                12'd315: toneL = `lg;
                12'd316: toneL = `lg;
                12'd317: toneL = `lg;
                12'd318: toneL = `lg;
                12'd319: toneL = `lg;
                12'd320: toneL = `la;
                12'd321: toneL = `la;
                12'd322: toneL = `la;
                12'd323: toneL = `la;
                12'd324: toneL = `la;
                12'd325: toneL = `la;
                12'd326: toneL = `la;
                12'd327: toneL = `la;
                12'd328: toneL = `la;
                12'd329: toneL = `la;
                12'd330: toneL = `la;
                12'd331: toneL = `la;
                12'd332: toneL = `la;
                12'd333: toneL = `la;
                12'd334: toneL = `la;
                12'd335: toneL = `la;
                12'd336: toneL = `la;
                12'd337: toneL = `la;
                12'd338: toneL = `la;
                12'd339: toneL = `la;
                12'd340: toneL = `la;
                12'd341: toneL = `la;
                12'd342: toneL = `la;
                12'd343: toneL = `la;
                12'd344: toneL = `la;
                12'd345: toneL = `la;
                12'd346: toneL = `la;
                12'd347: toneL = `la;
                12'd348: toneL = `la;
                12'd349: toneL = `la;
                12'd350: toneL = `la;
                12'd351: toneL = `la;
                12'd352: toneL = `la;
                12'd353: toneL = `la;
                12'd354: toneL = `la;
                12'd355: toneL = `la;
                12'd356: toneL = `la;
                12'd357: toneL = `la;
                12'd358: toneL = `la;
                12'd359: toneL = `la;
                12'd360: toneL = `la;
                12'd361: toneL = `la;
                12'd362: toneL = `la;
                12'd363: toneL = `la;
                12'd364: toneL = `la;
                12'd365: toneL = `la;
                12'd366: toneL = `la;
                12'd367: toneL = `la;
                12'd368: toneL = `la;
                12'd369: toneL = `la;
                12'd370: toneL = `la;
                12'd371: toneL = `la;
                12'd372: toneL = `la;
                12'd373: toneL = `la;
                12'd374: toneL = `la;
                12'd375: toneL = `la;
                12'd376: toneL = `la;
                12'd377: toneL = `la;
                12'd378: toneL = `la;
                12'd379: toneL = `la;
                12'd380: toneL = `la;
                12'd381: toneL = `la;
                12'd382: toneL = `la;
                12'd383: toneL = `la;
                12'd384: toneL = `g;
                12'd385: toneL = `g;
                12'd386: toneL = `g;
                12'd387: toneL = `g;
                12'd388: toneL = `g;
                12'd389: toneL = `g;
                12'd390: toneL = `g;
                12'd391: toneL = `g;
                12'd392: toneL = `g;
                12'd393: toneL = `g;
                12'd394: toneL = `g;
                12'd395: toneL = `g;
                12'd396: toneL = `g;
                12'd397: toneL = `g;
                12'd398: toneL = `g;
                12'd399: toneL = `sil;
                12'd400: toneL = `g;
                12'd401: toneL = `g;
                12'd402: toneL = `g;
                12'd403: toneL = `g;
                12'd404: toneL = `g;
                12'd405: toneL = `g;
                12'd406: toneL = `g;
                12'd407: toneL = `g;
                12'd408: toneL = `sf;
                12'd409: toneL = `sf;
                12'd410: toneL = `sf;
                12'd411: toneL = `sf;
                12'd412: toneL = `g;
                12'd413: toneL = `g;
                12'd414: toneL = `g;
                12'd415: toneL = `g;
                12'd416: toneL = `g;
                12'd417: toneL = `g;
                12'd418: toneL = `g;
                12'd419: toneL = `g;
                12'd420: toneL = `g;
                12'd421: toneL = `g;
                12'd422: toneL = `g;
                12'd423: toneL = `g;
                12'd424: toneL = `g;
                12'd425: toneL = `g;
                12'd426: toneL = `g;
                12'd427: toneL = `g;
                12'd428: toneL = `sil;
                12'd429: toneL = `sil;
                12'd430: toneL = `sil;
                12'd431: toneL = `sil;
                12'd432: toneL = `sil;
                12'd433: toneL = `sil;
                12'd434: toneL = `sil;
                12'd435: toneL = `sil;
                12'd436: toneL = `sil;
                12'd437: toneL = `sil;
                12'd438: toneL = `sil;
                12'd439: toneL = `sil;
                12'd440: toneL = `sil;
                12'd441: toneL = `sil;
                12'd442: toneL = `sil;
                12'd443: toneL = `sil;
                12'd444: toneL = `sil;
                12'd445: toneL = `sil;
                12'd446: toneL = `sil;
                12'd447: toneL = `sil;
                12'd448: toneL = `sil;
                12'd449: toneL = `sil;
                12'd450: toneL = `sil;
                12'd451: toneL = `sil;
                12'd452: toneL = `sil;
                12'd453: toneL = `sil;
                12'd454: toneL = `sil;
                12'd455: toneL = `sil;
                12'd456: toneL = `sil;
                12'd457: toneL = `sil;
                12'd458: toneL = `sil;
                12'd459: toneL = `sil;
                12'd460: toneL = `sil;
                12'd461: toneL = `sil;
                12'd462: toneL = `sil;
                12'd463: toneL = `sil;
                12'd464: toneL = `sil;
                12'd465: toneL = `sil;
                12'd466: toneL = `sil;
                12'd467: toneL = `sil;
                12'd468: toneL = `sil;
                12'd469: toneL = `sil;
                12'd470: toneL = `sil;
                12'd471: toneL = `sil;
                12'd472: toneL = `sil;
                12'd473: toneL = `sil;
                12'd474: toneL = `sil;
                12'd475: toneL = `sil;
                12'd476: toneL = `sil;
                12'd477: toneL = `sil;
                12'd478: toneL = `sil;
                12'd479: toneL = `sil;
                12'd480: toneL = `sil;
                12'd481: toneL = `sil;
                12'd482: toneL = `sil;
                12'd483: toneL = `sil;
                12'd484: toneL = `sil;
                12'd485: toneL = `sil;
                12'd486: toneL = `sil;
                12'd487: toneL = `sil;
                12'd488: toneL = `d;
                12'd489: toneL = `d;
                12'd490: toneL = `d;
                12'd491: toneL = `d;
                12'd492: toneL = `d;
                12'd493: toneL = `d;
                12'd494: toneL = `d;
                12'd495: toneL = `d;
                12'd496: toneL = `c;
                12'd497: toneL = `c;
                12'd498: toneL = `c;
                12'd499: toneL = `c;
                12'd500: toneL = `c;
                12'd501: toneL = `c;
                12'd502: toneL = `c;
                12'd503: toneL = `c;
                12'd504: toneL = `lg;
                12'd505: toneL = `lg;
                12'd506: toneL = `lg;
                12'd507: toneL = `lg;
                12'd508: toneL = `lg;
                12'd509: toneL = `lg;
                12'd510: toneL = `lg;
                12'd511: toneL = `lg;
                12'd512: toneL = `sil;
                12'd513: toneL = `sil;
                12'd514: toneL = `sil;
                12'd515: toneL = `sil;
                12'd516: toneL = `sil;
                12'd517: toneL = `sil;
                12'd518: toneL = `sil;
                12'd519: toneL = `sil;
                12'd520: toneL = `c;
                12'd521: toneL = `c;
                12'd522: toneL = `c;
                12'd523: toneL = `c;
                12'd524: toneL = `c;
                12'd525: toneL = `c;
                12'd526: toneL = `c;
                12'd527: toneL = `c;
                12'd528: toneL = `d;
                12'd529: toneL = `d;
                12'd530: toneL = `d;
                12'd531: toneL = `d;
                12'd532: toneL = `d;
                12'd533: toneL = `d;
                12'd534: toneL = `d;
                12'd535: toneL = `d;
                12'd536: toneL = `e;
                12'd537: toneL = `e;
                12'd538: toneL = `e;
                12'd539: toneL = `e;
                12'd540: toneL = `e;
                12'd541: toneL = `e;
                12'd542: toneL = `e;
                12'd543: toneL = `e;
                12'd544: toneL = `sil;
                12'd545: toneL = `sil;
                12'd546: toneL = `sil;
                12'd547: toneL = `sil;
                12'd548: toneL = `sil;
                12'd549: toneL = `sil;
                12'd550: toneL = `sil;
                12'd551: toneL = `sil;
                12'd552: toneL = `lg;
                12'd553: toneL = `lg;
                12'd554: toneL = `lg;
                12'd555: toneL = `lg;
                12'd556: toneL = `lg;
                12'd557: toneL = `lg;
                12'd558: toneL = `lg;
                12'd559: toneL = `lg;
                12'd560: toneL = `lg;
                12'd561: toneL = `lg;
                12'd562: toneL = `lg;
                12'd563: toneL = `lg;
                12'd564: toneL = `lg;
                12'd565: toneL = `lg;
                12'd566: toneL = `lg;
                12'd567: toneL = `lg;
                12'd568: toneL = `la;
                12'd569: toneL = `la;
                12'd570: toneL = `la;
                12'd571: toneL = `la;
                12'd572: toneL = `la;
                12'd573: toneL = `la;
                12'd574: toneL = `la;
                12'd575: toneL = `la;
                12'd576: toneL = `sil;
                12'd577: toneL = `sil;
                12'd578: toneL = `sil;
                12'd579: toneL = `sil;
                12'd580: toneL = `sil;
                12'd581: toneL = `sil;
                12'd582: toneL = `sil;
                12'd583: toneL = `sil;
                12'd584: toneL = `sil;
                12'd585: toneL = `sil;
                12'd586: toneL = `sil;
                12'd587: toneL = `sil;
                12'd588: toneL = `sil;
                12'd589: toneL = `sil;
                12'd590: toneL = `sil;
                12'd591: toneL = `sil;
                12'd592: toneL = `sil;
                12'd593: toneL = `sil;
                12'd594: toneL = `sil;
                12'd595: toneL = `sil;
                12'd596: toneL = `sil;
                12'd597: toneL = `sil;
                12'd598: toneL = `sil;
                12'd599: toneL = `sil;
                12'd600: toneL = `sil;
                12'd601: toneL = `sil;
                12'd602: toneL = `sil;
                12'd603: toneL = `sil;
                12'd604: toneL = `sil;
                12'd605: toneL = `sil;
                12'd606: toneL = `sil;
                12'd607: toneL = `sil;
                12'd608: toneL = `lb;
                12'd609: toneL = `lb;
                12'd610: toneL = `lb;
                12'd611: toneL = `lb;
                12'd612: toneL = `lb;
                12'd613: toneL = `lb;
                12'd614: toneL = `lb;
                12'd615: toneL = `lb;
                12'd616: toneL = `lb;
                12'd617: toneL = `lb;
                12'd618: toneL = `lb;
                12'd619: toneL = `lb;
                12'd620: toneL = `lb;
                12'd621: toneL = `lb;
                12'd622: toneL = `lb;
                12'd623: toneL = `lb;
                12'd624: toneL = `lf;
                12'd625: toneL = `lf;
                12'd626: toneL = `lf;
                12'd627: toneL = `lf;
                12'd628: toneL = `lf;
                12'd629: toneL = `lf;
                12'd630: toneL = `lf;
                12'd631: toneL = `lf;
                12'd632: toneL = `lf;
                12'd633: toneL = `lf;
                12'd634: toneL = `lf;
                12'd635: toneL = `lf;
                12'd636: toneL = `lf;
                12'd637: toneL = `lf;
                12'd638: toneL = `lf;
                12'd639: toneL = `lf;
                12'd640: toneL = `llb;
                12'd641: toneL = `llb;
                12'd642: toneL = `llb;
                12'd643: toneL = `llb;
                12'd644: toneL = `llb;
                12'd645: toneL = `llb;
                12'd646: toneL = `llb;
                12'd647: toneL = `llb;
                12'd648: toneL = `llb;
                12'd649: toneL = `llb;
                12'd650: toneL = `llb;
                12'd651: toneL = `llb;
                12'd652: toneL = `llb;
                12'd653: toneL = `llb;
                12'd654: toneL = `llb;
                12'd655: toneL = `llb;
                12'd656: toneL = `lg;
                12'd657: toneL = `lg;
                12'd658: toneL = `lg;
                12'd659: toneL = `lg;
                12'd660: toneL = `lg;
                12'd661: toneL = `lg;
                12'd662: toneL = `lg;
                12'd663: toneL = `lg;
                12'd664: toneL = `lg;
                12'd665: toneL = `lg;
                12'd666: toneL = `lg;
                12'd667: toneL = `lg;
                12'd668: toneL = `lg;
                12'd669: toneL = `lg;
                12'd670: toneL = `lg;
                12'd671: toneL = `lg;
                12'd672: toneL = `e;
                12'd673: toneL = `e;
                12'd674: toneL = `e;
                12'd675: toneL = `e;
                12'd676: toneL = `e;
                12'd677: toneL = `e;
                12'd678: toneL = `e;
                12'd679: toneL = `e;
                12'd680: toneL = `e;
                12'd681: toneL = `e;
                12'd682: toneL = `e;
                12'd683: toneL = `e;
                12'd684: toneL = `e;
                12'd685: toneL = `e;
                12'd686: toneL = `e;
                12'd687: toneL = `e;
                12'd688: toneL = `e;
                12'd689: toneL = `e;
                12'd690: toneL = `e;
                12'd691: toneL = `e;
                12'd692: toneL = `e;
                12'd693: toneL = `e;
                12'd694: toneL = `e;
                12'd695: toneL = `e;
                12'd696: toneL = `e;
                12'd697: toneL = `e;
                12'd698: toneL = `e;
                12'd699: toneL = `e;
                12'd700: toneL = `e;
                12'd701: toneL = `e;
                12'd702: toneL = `e;
                12'd703: toneL = `e;
                12'd704: toneL = `sil;
                12'd705: toneL = `sil;
                12'd706: toneL = `sil;
                12'd707: toneL = `sil;
                12'd708: toneL = `sil;
                12'd709: toneL = `sil;
                12'd710: toneL = `sil;
                12'd711: toneL = `sil;
                12'd712: toneL = `sil;
                12'd713: toneL = `sil;
                12'd714: toneL = `sil;
                12'd715: toneL = `sil;
                12'd716: toneL = `sil;
                12'd717: toneL = `sil;
                12'd718: toneL = `sil;
                12'd719: toneL = `sil;
                12'd720: toneL = `sil;
                12'd721: toneL = `sil;
                12'd722: toneL = `sil;
                12'd723: toneL = `sil;
                12'd724: toneL = `sil;
                12'd725: toneL = `sil;
                12'd726: toneL = `sil;
                12'd727: toneL = `sil;
                12'd728: toneL = `sil;
                12'd729: toneL = `sil;
                12'd730: toneL = `sil;
                12'd731: toneL = `sil;
                12'd732: toneL = `sil;
                12'd733: toneL = `sil;
                12'd734: toneL = `sil;
                12'd735: toneL = `sil;
                12'd736: toneL = `sil;
                12'd737: toneL = `sil;
                12'd738: toneL = `sil;
                12'd739: toneL = `sil;
                12'd740: toneL = `sil;
                12'd741: toneL = `sil;
                12'd742: toneL = `sil;
                12'd743: toneL = `sil;
                12'd744: toneL = `c;
                12'd745: toneL = `c;
                12'd746: toneL = `c;
                12'd747: toneL = `c;
                12'd748: toneL = `c;
                12'd749: toneL = `c;
                12'd750: toneL = `c;
                12'd751: toneL = `c;
                12'd752: toneL = `d;
                12'd753: toneL = `d;
                12'd754: toneL = `d;
                12'd755: toneL = `d;
                12'd756: toneL = `d;
                12'd757: toneL = `d;
                12'd758: toneL = `d;
                12'd759: toneL = `d;
                12'd760: toneL = `e;
                12'd761: toneL = `e;
                12'd762: toneL = `e;
                12'd763: toneL = `e;
                12'd764: toneL = `e;
                12'd765: toneL = `e;
                12'd766: toneL = `e;
                12'd767: toneL = `e;
                12'd768: toneL = `sil;
                12'd769: toneL = `sil;
                12'd770: toneL = `sil;
                12'd771: toneL = `sil;
                12'd772: toneL = `sil;
                12'd773: toneL = `sil;
                12'd774: toneL = `sil;
                12'd775: toneL = `sil;
                12'd776: toneL = `lg;
                12'd777: toneL = `lg;
                12'd778: toneL = `lg;
                12'd779: toneL = `lg;
                12'd780: toneL = `lg;
                12'd781: toneL = `lg;
                12'd782: toneL = `lg;
                12'd783: toneL = `lg;
                12'd784: toneL = `lg;
                12'd785: toneL = `lg;
                12'd786: toneL = `lg;
                12'd787: toneL = `lg;
                12'd788: toneL = `lg;
                12'd789: toneL = `lg;
                12'd790: toneL = `lg;
                12'd791: toneL = `lg;
                12'd792: toneL = `la;
                12'd793: toneL = `la;
                12'd794: toneL = `la;
                12'd795: toneL = `la;
                12'd796: toneL = `la;
                12'd797: toneL = `la;
                12'd798: toneL = `la;
                12'd799: toneL = `la;
                12'd800: toneL = `la;
                12'd801: toneL = `la;
                12'd802: toneL = `la;
                12'd803: toneL = `la;
                12'd804: toneL = `la;
                12'd805: toneL = `la;
                12'd806: toneL = `la;
                12'd807: toneL = `la;
                12'd808: toneL = `la;
                12'd809: toneL = `la;
                12'd810: toneL = `la;
                12'd811: toneL = `la;
                12'd812: toneL = `la;
                12'd813: toneL = `la;
                12'd814: toneL = `la;
                12'd815: toneL = `la;
                12'd816: toneL = `la;
                12'd817: toneL = `la;
                12'd818: toneL = `la;
                12'd819: toneL = `la;
                12'd820: toneL = `la;
                12'd821: toneL = `la;
                12'd822: toneL = `la;
                12'd823: toneL = `la;
                12'd824: toneL = `sil;
                12'd825: toneL = `sil;
                12'd826: toneL = `sil;
                12'd827: toneL = `sil;
                12'd828: toneL = `sil;
                12'd829: toneL = `sil;
                12'd830: toneL = `sil;
                12'd831: toneL = `sil;
                12'd832: toneL = `d;
                12'd833: toneL = `d;
                12'd834: toneL = `d;
                12'd835: toneL = `d;
                12'd836: toneL = `d;
                12'd837: toneL = `d;
                12'd838: toneL = `d;
                12'd839: toneL = `d;
                12'd840: toneL = `d;
                12'd841: toneL = `d;
                12'd842: toneL = `d;
                12'd843: toneL = `d;
                12'd844: toneL = `d;
                12'd845: toneL = `d;
                12'd846: toneL = `d;
                12'd847: toneL = `d;
                12'd848: toneL = `sf;
                12'd849: toneL = `sf;
                12'd850: toneL = `sf;
                12'd851: toneL = `sf;
                12'd852: toneL = `sf;
                12'd853: toneL = `sf;
                12'd854: toneL = `sf;
                12'd855: toneL = `sf;
                12'd856: toneL = `sf;
                12'd857: toneL = `sf;
                12'd858: toneL = `sf;
                12'd859: toneL = `sf;
                12'd860: toneL = `sf;
                12'd861: toneL = `sf;
                12'd862: toneL = `sf;
                12'd863: toneL = `sf;
                12'd864: toneL = `sil;
                12'd865: toneL = `sil;
                12'd866: toneL = `sil;
                12'd867: toneL = `sil;
                12'd868: toneL = `sil;
                12'd869: toneL = `sil;
                12'd870: toneL = `sil;
                12'd871: toneL = `sil;
                12'd872: toneL = `e;
                12'd873: toneL = `e;
                12'd874: toneL = `e;
                12'd875: toneL = `e;
                12'd876: toneL = `e;
                12'd877: toneL = `e;
                12'd878: toneL = `e;
                12'd879: toneL = `e;
                12'd880: toneL = `e;
                12'd881: toneL = `e;
                12'd882: toneL = `e;
                12'd883: toneL = `e;
                12'd884: toneL = `e;
                12'd885: toneL = `e;
                12'd886: toneL = `e;
                12'd887: toneL = `e;
                12'd888: toneL = `sil;
                12'd889: toneL = `sil;
                12'd890: toneL = `sil;
                12'd891: toneL = `sil;
                12'd892: toneL = `sil;
                12'd893: toneL = `sil;
                12'd894: toneL = `sil;
                12'd895: toneL = `sil;
                12'd896: toneL = `sil;
                12'd897: toneL = `sil;
                12'd898: toneL = `sil;
                12'd899: toneL = `sil;
                12'd900: toneL = `sil;
                12'd901: toneL = `sil;
                12'd902: toneL = `sil;
                12'd903: toneL = `sil;
                12'd904: toneL = `sil;
                12'd905: toneL = `sil;
                12'd906: toneL = `sil;
                12'd907: toneL = `sil;
                12'd908: toneL = `sil;
                12'd909: toneL = `sil;
                12'd910: toneL = `sil;
                12'd911: toneL = `sil;
                12'd912: toneL = `sil;
                12'd913: toneL = `sil;
                12'd914: toneL = `sil;
                12'd915: toneL = `sil;
                12'd916: toneL = `sil;
                12'd917: toneL = `sil;
                12'd918: toneL = `sil;
                12'd919: toneL = `sil;
                12'd920: toneL = `c;
                12'd921: toneL = `c;
                12'd922: toneL = `c;
                12'd923: toneL = `c;
                12'd924: toneL = `c;
                12'd925: toneL = `c;
                12'd926: toneL = `c;
                12'd927: toneL = `c;
                12'd928: toneL = `c;
                12'd929: toneL = `c;
                12'd930: toneL = `c;
                12'd931: toneL = `c;
                12'd932: toneL = `c;
                12'd933: toneL = `c;
                12'd934: toneL = `c;
                12'd935: toneL = `c;
                12'd936: toneL = `c;
                12'd937: toneL = `c;
                12'd938: toneL = `c;
                12'd939: toneL = `c;
                12'd940: toneL = `c;
                12'd941: toneL = `c;
                12'd942: toneL = `c;
                12'd943: toneL = `c;
                12'd944: toneL = `c;
                12'd945: toneL = `c;
                12'd946: toneL = `c;
                12'd947: toneL = `c;
                12'd948: toneL = `c;
                12'd949: toneL = `c;
                12'd950: toneL = `c;
                12'd951: toneL = `c;
                12'd952: toneL = `sil;
                12'd953: toneL = `sil;
                12'd954: toneL = `sil;
                12'd955: toneL = `sil;
                12'd956: toneL = `sil;
                12'd957: toneL = `sil;
                12'd958: toneL = `sil;
                12'd959: toneL = `sil;
                12'd960: toneL = `c;
                12'd961: toneL = `c;
                12'd962: toneL = `c;
                12'd963: toneL = `c;
                12'd964: toneL = `c;
                12'd965: toneL = `c;
                12'd966: toneL = `c;
                12'd967: toneL = `c;
                12'd968: toneL = `lb;
                12'd969: toneL = `lb;
                12'd970: toneL = `lb;
                12'd971: toneL = `lb;
                12'd972: toneL = `lb;
                12'd973: toneL = `lb;
                12'd974: toneL = `lb;
                12'd975: toneL = `lb;
                12'd976: toneL = `lsa;
                12'd977: toneL = `lsa;
                12'd978: toneL = `lsa;
                12'd979: toneL = `lsa;
                12'd980: toneL = `lsa;
                12'd981: toneL = `lsa;
                12'd982: toneL = `lsa;
                12'd983: toneL = `lsa;
                12'd984: toneL = `lsa;
                12'd985: toneL = `lsa;
                12'd986: toneL = `lsa;
                12'd987: toneL = `lsa;
                12'd988: toneL = `lsa;
                12'd989: toneL = `lsa;
                12'd990: toneL = `lsa;
                12'd991: toneL = `lsa;
                12'd992: toneL = `sil;
                12'd993: toneL = `sil;
                12'd994: toneL = `sil;
                12'd995: toneL = `sil;
                12'd996: toneL = `sil;
                12'd997: toneL = `sil;
                12'd998: toneL = `sil;
                12'd999: toneL = `sil;
                12'd1000: toneL = `sil;
                12'd1001: toneL = `sil;
                12'd1002: toneL = `sil;
                12'd1003: toneL = `sil;
                12'd1004: toneL = `sil;
                12'd1005: toneL = `sil;
                12'd1006: toneL = `sil;
                12'd1007: toneL = `sil;
                12'd1008: toneL = `la;
                12'd1009: toneL = `la;
                12'd1010: toneL = `la;
                12'd1011: toneL = `la;
                12'd1012: toneL = `la;
                12'd1013: toneL = `la;
                12'd1014: toneL = `la;
                12'd1015: toneL = `la;
                12'd1016: toneL = `lb;
                12'd1017: toneL = `lb;
                12'd1018: toneL = `lb;
                12'd1019: toneL = `lb;
                12'd1020: toneL = `lb;
                12'd1021: toneL = `lb;
                12'd1022: toneL = `lb;
                12'd1023: toneL = `lb;
                12'd1024: toneL = `c;
                12'd1025: toneL = `c;
                12'd1026: toneL = `c;
                12'd1027: toneL = `c;
                12'd1028: toneL = `c;
                12'd1029: toneL = `c;
                12'd1030: toneL = `c;
                12'd1031: toneL = `c;
                12'd1032: toneL = `d;
                12'd1033: toneL = `d;
                12'd1034: toneL = `d;
                12'd1035: toneL = `d;
                12'd1036: toneL = `d;
                12'd1037: toneL = `d;
                12'd1038: toneL = `d;
                12'd1039: toneL = `d;
                12'd1040: toneL = `f;
                12'd1041: toneL = `f;
                12'd1042: toneL = `f;
                12'd1043: toneL = `f;
                12'd1044: toneL = `f;
                12'd1045: toneL = `f;
                12'd1046: toneL = `f;
                12'd1047: toneL = `f;
                12'd1048: toneL = `d;
                12'd1049: toneL = `d;
                12'd1050: toneL = `d;
                12'd1051: toneL = `d;
                12'd1052: toneL = `d;
                12'd1053: toneL = `d;
                12'd1054: toneL = `d;
                12'd1055: toneL = `d;
                12'd1056: toneL = `c;
                12'd1057: toneL = `c;
                12'd1058: toneL = `c;
                12'd1059: toneL = `c;
                12'd1060: toneL = `c;
                12'd1061: toneL = `c;
                12'd1062: toneL = `c;
                12'd1063: toneL = `c;
                12'd1064: toneL = `c;
                12'd1065: toneL = `c;
                12'd1066: toneL = `c;
                12'd1067: toneL = `c;
                12'd1068: toneL = `c;
                12'd1069: toneL = `c;
                12'd1070: toneL = `c;
                12'd1071: toneL = `c;
                12'd1072: toneL = `lg;
                12'd1073: toneL = `lg;
                12'd1074: toneL = `lg;
                12'd1075: toneL = `lg;
                12'd1076: toneL = `lg;
                12'd1077: toneL = `lg;
                12'd1078: toneL = `lg;
                12'd1079: toneL = `lg;
                12'd1080: toneL = `lg;
                12'd1081: toneL = `lg;
                12'd1082: toneL = `lg;
                12'd1083: toneL = `lg;
                12'd1084: toneL = `lg;
                12'd1085: toneL = `lg;
                12'd1086: toneL = `lg;
                12'd1087: toneL = `lg;
                12'd1088: toneL = `sil;
                12'd1089: toneL = `sil;
                12'd1090: toneL = `sil;
                12'd1091: toneL = `sil;
                12'd1092: toneL = `sil;
                12'd1093: toneL = `sil;
                12'd1094: toneL = `sil;
                12'd1095: toneL = `sil;
                12'd1096: toneL = `c;
                12'd1097: toneL = `c;
                12'd1098: toneL = `c;
                12'd1099: toneL = `c;
                12'd1100: toneL = `c;
                12'd1101: toneL = `c;
                12'd1102: toneL = `c;
                12'd1103: toneL = `c;
                12'd1104: toneL = `lb;
                12'd1105: toneL = `lb;
                12'd1106: toneL = `lb;
                12'd1107: toneL = `lb;
                12'd1108: toneL = `lb;
                12'd1109: toneL = `lb;
                12'd1110: toneL = `lb;
                12'd1111: toneL = `lb;
                12'd1112: toneL = `sil;
                12'd1113: toneL = `sil;
                12'd1114: toneL = `sil;
                12'd1115: toneL = `sil;
                12'd1116: toneL = `sil;
                12'd1117: toneL = `sil;
                12'd1118: toneL = `sil;
                12'd1119: toneL = `sil;
                12'd1120: toneL = `sil;
                12'd1121: toneL = `sil;
                12'd1122: toneL = `sil;
                12'd1123: toneL = `sil;
                12'd1124: toneL = `sil;
                12'd1125: toneL = `sil;
                12'd1126: toneL = `sil;
                12'd1127: toneL = `sil;
                12'd1128: toneL = `sil;
                12'd1129: toneL = `sil;
                12'd1130: toneL = `sil;
                12'd1131: toneL = `sil;
                12'd1132: toneL = `sil;
                12'd1133: toneL = `sil;
                12'd1134: toneL = `sil;
                12'd1135: toneL = `sil;
                12'd1136: toneL = `sil;
                12'd1137: toneL = `sil;
                12'd1138: toneL = `sil;
                12'd1139: toneL = `sil;
                12'd1140: toneL = `sil;
                12'd1141: toneL = `sil;
                12'd1142: toneL = `sil;
                12'd1143: toneL = `sil;
                12'd1144: toneL = `sil;
                12'd1145: toneL = `sil;
                12'd1146: toneL = `sil;
                12'd1147: toneL = `sil;
                12'd1148: toneL = `sil;
                12'd1149: toneL = `sil;
                12'd1150: toneL = `sil;
                12'd1151: toneL = `sil;
                12'd1152: toneL = `a;
                12'd1153: toneL = `a;
                12'd1154: toneL = `a;
                12'd1155: toneL = `a;
                12'd1156: toneL = `a;
                12'd1157: toneL = `a;
                12'd1158: toneL = `a;
                12'd1159: toneL = `a;
                12'd1160: toneL = `b;
                12'd1161: toneL = `b;
                12'd1162: toneL = `b;
                12'd1163: toneL = `b;
                12'd1164: toneL = `b;
                12'd1165: toneL = `b;
                12'd1166: toneL = `b;
                12'd1167: toneL = `b;
                12'd1168: toneL = `hc;
                12'd1169: toneL = `hc;
                12'd1170: toneL = `hc;
                12'd1171: toneL = `hc;
                12'd1172: toneL = `hc;
                12'd1173: toneL = `hc;
                12'd1174: toneL = `hc;
                12'd1175: toneL = `hc;
                12'd1176: toneL = `b;
                12'd1177: toneL = `b;
                12'd1178: toneL = `b;
                12'd1179: toneL = `b;
                12'd1180: toneL = `b;
                12'd1181: toneL = `b;
                12'd1182: toneL = `b;
                12'd1183: toneL = `b;
                12'd1184: toneL = `a;
                12'd1185: toneL = `a;
                12'd1186: toneL = `a;
                12'd1187: toneL = `a;
                12'd1188: toneL = `a;
                12'd1189: toneL = `a;
                12'd1190: toneL = `a;
                12'd1191: toneL = `a;
                12'd1192: toneL = `a;
                12'd1193: toneL = `a;
                12'd1194: toneL = `a;
                12'd1195: toneL = `a;
                12'd1196: toneL = `a;
                12'd1197: toneL = `a;
                12'd1198: toneL = `a;
                12'd1199: toneL = `a;
                12'd1200: toneL = `e;
                12'd1201: toneL = `e;
                12'd1202: toneL = `e;
                12'd1203: toneL = `e;
                12'd1204: toneL = `e;
                12'd1205: toneL = `e;
                12'd1206: toneL = `e;
                12'd1207: toneL = `e;
                12'd1208: toneL = `e;
                12'd1209: toneL = `e;
                12'd1210: toneL = `e;
                12'd1211: toneL = `e;
                12'd1212: toneL = `e;
                12'd1213: toneL = `e;
                12'd1214: toneL = `e;
                12'd1215: toneL = `e;
                12'd1216: toneL = `c;
                12'd1217: toneL = `c;
                12'd1218: toneL = `c;
                12'd1219: toneL = `c;
                12'd1220: toneL = `c;
                12'd1221: toneL = `c;
                12'd1222: toneL = `c;
                12'd1223: toneL = `c;
                12'd1224: toneL = `hc;
                12'd1225: toneL = `hc;
                12'd1226: toneL = `hc;
                12'd1227: toneL = `hc;
                12'd1228: toneL = `hc;
                12'd1229: toneL = `hc;
                12'd1230: toneL = `hc;
                12'd1231: toneL = `hc;
                12'd1232: toneL = `sil;
                12'd1233: toneL = `sil;
                12'd1234: toneL = `sil;
                12'd1235: toneL = `sil;
                12'd1236: toneL = `sil;
                12'd1237: toneL = `sil;
                12'd1238: toneL = `sil;
                12'd1239: toneL = `sil;
                12'd1240: toneL = `sil;
                12'd1241: toneL = `sil;
                12'd1242: toneL = `sil;
                12'd1243: toneL = `sil;
                12'd1244: toneL = `sil;
                12'd1245: toneL = `sil;
                12'd1246: toneL = `sil;
                12'd1247: toneL = `sil;
                12'd1248: toneL = `sil;
                12'd1249: toneL = `sil;
                12'd1250: toneL = `sil;
                12'd1251: toneL = `sil;
                12'd1252: toneL = `sil;
                12'd1253: toneL = `sil;
                12'd1254: toneL = `sil;
                12'd1255: toneL = `sil;
                12'd1256: toneL = `sil;
                12'd1257: toneL = `sil;
                12'd1258: toneL = `sil;
                12'd1259: toneL = `sil;
                12'd1260: toneL = `sil;
                12'd1261: toneL = `sil;
                12'd1262: toneL = `sil;
                12'd1263: toneL = `sil;
                12'd1264: toneL = `c;
                12'd1265: toneL = `c;
                12'd1266: toneL = `c;
                12'd1267: toneL = `c;
                12'd1268: toneL = `c;
                12'd1269: toneL = `c;
                12'd1270: toneL = `c;
                12'd1271: toneL = `c;
                12'd1272: toneL = `c;
                12'd1273: toneL = `c;
                12'd1274: toneL = `c;
                12'd1275: toneL = `c;
                12'd1276: toneL = `c;
                12'd1277: toneL = `c;
                12'd1278: toneL = `c;
                12'd1279: toneL = `sil;
                12'd1280: toneL = `c;
                12'd1281: toneL = `c;
                12'd1282: toneL = `c;
                12'd1283: toneL = `c;
                12'd1284: toneL = `c;
                12'd1285: toneL = `c;
                12'd1286: toneL = `c;
                12'd1287: toneL = `c;
                12'd1288: toneL = `c;
                12'd1289: toneL = `c;
                12'd1290: toneL = `c;
                12'd1291: toneL = `c;
                12'd1292: toneL = `c;
                12'd1293: toneL = `c;
                12'd1294: toneL = `c;
                12'd1295: toneL = `c;
                12'd1296: toneL = `lb;
                12'd1297: toneL = `lb;
                12'd1298: toneL = `lb;
                12'd1299: toneL = `lb;
                12'd1300: toneL = `lb;
                12'd1301: toneL = `lb;
                12'd1302: toneL = `lb;
                12'd1303: toneL = `lb;
                12'd1304: toneL = `lb;
                12'd1305: toneL = `lb;
                12'd1306: toneL = `lb;
                12'd1307: toneL = `lb;
                12'd1308: toneL = `lb;
                12'd1309: toneL = `lb;
                12'd1310: toneL = `lb;
                12'd1311: toneL = `lb;
                12'd1312: toneL = `c;
                12'd1313: toneL = `c;
                12'd1314: toneL = `c;
                12'd1315: toneL = `c;
                12'd1316: toneL = `c;
                12'd1317: toneL = `c;
                12'd1318: toneL = `c;
                12'd1319: toneL = `c;
                12'd1320: toneL = `lb;
                12'd1321: toneL = `lb;
                12'd1322: toneL = `lb;
                12'd1323: toneL = `lb;
                12'd1324: toneL = `lb;
                12'd1325: toneL = `lb;
                12'd1326: toneL = `lb;
                12'd1327: toneL = `lb;
                12'd1328: toneL = `la;
                12'd1329: toneL = `la;
                12'd1330: toneL = `la;
                12'd1331: toneL = `la;
                12'd1332: toneL = `la;
                12'd1333: toneL = `la;
                12'd1334: toneL = `la;
                12'd1335: toneL = `la;
                12'd1336: toneL = `lb;
                12'd1337: toneL = `lb;
                12'd1338: toneL = `lb;
                12'd1339: toneL = `lb;
                12'd1340: toneL = `lb;
                12'd1341: toneL = `lb;
                12'd1342: toneL = `lb;
                12'd1343: toneL = `lb;
                12'd1344: toneL = `c;
                12'd1345: toneL = `c;
                12'd1346: toneL = `c;
                12'd1347: toneL = `c;
                12'd1348: toneL = `c;
                12'd1349: toneL = `c;
                12'd1350: toneL = `c;
                12'd1351: toneL = `c;
                12'd1352: toneL = `g;
                12'd1353: toneL = `g;
                12'd1354: toneL = `g;
                12'd1355: toneL = `g;
                12'd1356: toneL = `g;
                12'd1357: toneL = `g;
                12'd1358: toneL = `g;
                12'd1359: toneL = `g;
                12'd1360: toneL = `sil;
                12'd1361: toneL = `sil;
                12'd1362: toneL = `sil;
                12'd1363: toneL = `sil;
                12'd1364: toneL = `sil;
                12'd1365: toneL = `sil;
                12'd1366: toneL = `sil;
                12'd1367: toneL = `sil;
                12'd1368: toneL = `sil;
                12'd1369: toneL = `sil;
                12'd1370: toneL = `sil;
                12'd1371: toneL = `sil;
                12'd1372: toneL = `sil;
                12'd1373: toneL = `sil;
                12'd1374: toneL = `sil;
                12'd1375: toneL = `sil;
                12'd1376: toneL = `b;
                12'd1377: toneL = `b;
                12'd1378: toneL = `b;
                12'd1379: toneL = `b;
                12'd1380: toneL = `b;
                12'd1381: toneL = `b;
                12'd1382: toneL = `b;
                12'd1383: toneL = `b;
                12'd1384: toneL = `b;
                12'd1385: toneL = `b;
                12'd1386: toneL = `b;
                12'd1387: toneL = `b;
                12'd1388: toneL = `b;
                12'd1389: toneL = `b;
                12'd1390: toneL = `b;
                12'd1391: toneL = `b;
                12'd1392: toneL = `b;
                12'd1393: toneL = `b;
                12'd1394: toneL = `b;
                12'd1395: toneL = `b;
                12'd1396: toneL = `b;
                12'd1397: toneL = `b;
                12'd1398: toneL = `b;
                12'd1399: toneL = `b;
                12'd1400: toneL = `b;
                12'd1401: toneL = `b;
                12'd1402: toneL = `b;
                12'd1403: toneL = `b;
                12'd1404: toneL = `b;
                12'd1405: toneL = `b;
                12'd1406: toneL = `b;
                12'd1407: toneL = `b;
                12'd1408: toneL = `f;
                12'd1409: toneL = `f;
                12'd1410: toneL = `f;
                12'd1411: toneL = `f;
                12'd1412: toneL = `f;
                12'd1413: toneL = `f;
                12'd1414: toneL = `f;
                12'd1415: toneL = `f;
                12'd1416: toneL = `lf;
                12'd1417: toneL = `lf;
                12'd1418: toneL = `lf;
                12'd1419: toneL = `lf;
                12'd1420: toneL = `lf;
                12'd1421: toneL = `lf;
                12'd1422: toneL = `lf;
                12'd1423: toneL = `lf;
                12'd1424: toneL = `g;
                12'd1425: toneL = `g;
                12'd1426: toneL = `g;
                12'd1427: toneL = `g;
                12'd1428: toneL = `g;
                12'd1429: toneL = `g;
                12'd1430: toneL = `g;
                12'd1431: toneL = `g;
                12'd1432: toneL = `lg;
                12'd1433: toneL = `lg;
                12'd1434: toneL = `lg;
                12'd1435: toneL = `lg;
                12'd1436: toneL = `lg;
                12'd1437: toneL = `lg;
                12'd1438: toneL = `lg;
                12'd1439: toneL = `lg;
                12'd1440: toneL = `b;
                12'd1441: toneL = `b;
                12'd1442: toneL = `b;
                12'd1443: toneL = `b;
                12'd1444: toneL = `b;
                12'd1445: toneL = `b;
                12'd1446: toneL = `b;
                12'd1447: toneL = `sil;
                12'd1448: toneL = `b;
                12'd1449: toneL = `b;
                12'd1450: toneL = `b;
                12'd1451: toneL = `b;
                12'd1452: toneL = `b;
                12'd1453: toneL = `b;
                12'd1454: toneL = `b;
                12'd1455: toneL = `b;
                12'd1456: toneL = `hc;
                12'd1457: toneL = `hc;
                12'd1458: toneL = `hc;
                12'd1459: toneL = `hc;
                12'd1460: toneL = `hc;
                12'd1461: toneL = `hc;
                12'd1462: toneL = `hc;
                12'd1463: toneL = `hc;
                12'd1464: toneL = `hc;
                12'd1465: toneL = `hc;
                12'd1466: toneL = `hc;
                12'd1467: toneL = `hc;
                12'd1468: toneL = `hc;
                12'd1469: toneL = `hc;
                12'd1470: toneL = `hc;
                12'd1471: toneL = `hc;
                12'd1472: toneL = `c;
                12'd1473: toneL = `c;
                12'd1474: toneL = `d;
                12'd1475: toneL = `d;
                12'd1476: toneL = `e;
                12'd1477: toneL = `e;
                12'd1478: toneL = `f;
                12'd1479: toneL = `f;
                12'd1480: toneL = `g;
                12'd1481: toneL = `g;
                12'd1482: toneL = `a;
                12'd1483: toneL = `a;
                12'd1484: toneL = `b;
                12'd1485: toneL = `b;
                12'd1486: toneL = `hc;
                12'd1487: toneL = `hc;
                12'd1488: toneL = `sil;
                12'd1489: toneL = `sil;
                12'd1490: toneL = `sil;
                12'd1491: toneL = `sil;
                12'd1492: toneL = `sil;
                12'd1493: toneL = `sil;
                12'd1494: toneL = `sil;
                12'd1495: toneL = `sil;
                12'd1496: toneL = `sil;
                12'd1497: toneL = `sil;
                12'd1498: toneL = `sil;
                12'd1499: toneL = `sil;
                12'd1500: toneL = `sil;
                12'd1501: toneL = `sil;
                12'd1502: toneL = `sil;
                12'd1503: toneL = `sil;
                12'd1504: toneL = `lllc;
                12'd1505: toneL = `lllc;
                12'd1506: toneL = `lllc;
                12'd1507: toneL = `lllc;
                12'd1508: toneL = `lllc;
                12'd1509: toneL = `lllc;
                12'd1510: toneL = `lllc;
                12'd1511: toneL = `lllc;
                12'd1512: toneL = `lllc;
                12'd1513: toneL = `lllc;
                12'd1514: toneL = `lllc;
                12'd1515: toneL = `lllc;
                12'd1516: toneL = `lllc;
                12'd1517: toneL = `lllc;
                12'd1518: toneL = `lllc;
                12'd1519: toneL = `lllc;
                12'd1520: toneL = `lllc;
                12'd1521: toneL = `lllc;
                12'd1522: toneL = `lllc;
                12'd1523: toneL = `lllc;
                12'd1524: toneL = `lllc;
                12'd1525: toneL = `lllc;
                12'd1526: toneL = `lllc;
                12'd1527: toneL = `lllc;
                12'd1528: toneL = `lllc;
                12'd1529: toneL = `lllc;
                12'd1530: toneL = `lllc;
                12'd1531: toneL = `lllc;
                12'd1532: toneL = `lllc;
                12'd1533: toneL = `lllc;
                12'd1534: toneL = `lllc;
                12'd1535: toneL = `lllc;
            default:toneL = `sil;
        endcase
    end
    else toneL = `sil;
end
endmodule